class c_1305_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1305_6;
    c_1305_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1111xz11zzz0xz1x101zx10z1xzz0x1xxzxzxxxxxzzzzzxxxxxxxxxxzxzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
