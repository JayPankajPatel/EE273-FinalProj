class c_320_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_320_6;
    c_320_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x10z1x0101xzx10z11010zxz1x1x001zxzxzzzzzzxxzxzzzxzzxzzxxxxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
