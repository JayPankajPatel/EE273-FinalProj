class c_1155_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1155_6;
    c_1155_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111x0x0z1z011zx10111zx1zzz001110xzzxxxzxxzxxzzzzzxzxzxzxxzzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
