class c_1790_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1790_6;
    c_1790_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01x1z0x1xx1x10zxx0zzz010xz00z1xxxxxxzzzzxzzxzzzxxxzzzzzxzzzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
