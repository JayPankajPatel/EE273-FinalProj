class c_1247_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1247_6;
    c_1247_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x10z00z000xx0xz0z0101xzzx0011x1zzxxxxzzzzzzzxzxzzxxzzxzxxxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
