class c_1806_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1806_6;
    c_1806_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z11z1zx0zx1xz10x00101zzzx1x1xzxzxxxxzxxzzxxxxxzxzxxzxxzzxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
