class c_1840_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1840_6;
    c_1840_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz011z10xx10xzx0z110zz101x00xz0zzzxxzzxzzzzzzxxxxzxzxzxzxxzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
