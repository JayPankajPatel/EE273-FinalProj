class c_1565_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1565_6;
    c_1565_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz1zx0x0010100xzx0z0zzxxx10xz000zxxzxxzzxzzzzxzzzzzzzxzzxzzxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
