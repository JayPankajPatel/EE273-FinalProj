class c_486_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_486_6;
    c_486_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00x10x0xz1zz0z0xz00xxxzz010xxzzxxxzxzxzxxzzxxxzxzzzzzxzzzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
