class c_1546_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1546_6;
    c_1546_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzx010z0x100x1zxx0x0x1zx1xz10zz0xxzxxzxzxxzxzzzxzxzxxxzzzzzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
