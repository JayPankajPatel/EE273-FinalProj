class c_1784_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1784_6;
    c_1784_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zx1x1z101zxx1zxzxxzx0xxzx0zzz1zxzxzxxxxzxzxzzxxxxxxxxxzxzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
