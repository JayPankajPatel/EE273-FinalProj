class c_1628_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1628_6;
    c_1628_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx1zx1z1111z1x0x0xx0x1z000zxx101zzxxxxzxxxzzxxxxxxxzzzxzzxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
