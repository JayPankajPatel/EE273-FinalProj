class c_532_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_532_6;
    c_532_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx1xxx1zxz1zz00x100x0zxxz0zzx110xxzxzzzxxzzzxxxxxxzzxxzzzxxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
