class c_1814_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1814_6;
    c_1814_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x00xzzx11xz100100x1zz01xzz001z0xxzxxzzzzxxzzzxzxxzxzzxzxzzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
