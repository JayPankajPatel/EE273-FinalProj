class c_1058_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1058_6;
    c_1058_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x000zz1zx1xzz1z0x1xz1z01z0z0xzzxzxxxxxzxxzxzzxzzxxzxxzzzzxzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
