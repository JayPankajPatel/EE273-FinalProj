class c_1485_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1485_6;
    c_1485_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0zxx0x00z01x1zx1x0xzxx11z0xx0xzzxxzxxxxxzxzzzxzxzzxxxxzzxxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
