class c_1373_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1373_6;
    c_1373_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10010z0011x1xxz0z0x01xxxxzzz1z0zxzxzzxzzzzzzxxxxzxzxzxxzzzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
