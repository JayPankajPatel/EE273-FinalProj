class c_1542_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1542_6;
    c_1542_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "010zx0x01xxzxxxx0x1zz0001100x1z1zzxzxxzxzxzxxxzxxzzxxzxzxzxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
