class c_908_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_908_6;
    c_908_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz1x0xzz10x0z1xz01zxxzzz0zx0zx1xzxxxzzxxxxzzzxzzxzzxxzxxzzzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
