class c_1314_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1314_6;
    c_1314_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01100xz11xz10z011xzx1zx0xz00z1x0xzxzxzzzxxzxzzzzxzxzxzxzzzzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
