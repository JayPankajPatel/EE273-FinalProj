class c_1379_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1379_6;
    c_1379_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx1zz1z10z0zx1z0zxzxzx10101z10x1xxzxxxxxzzxzzzzzxxzzzzxzxzzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
