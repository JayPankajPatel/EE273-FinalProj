class c_731_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_731_6;
    c_731_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x1z11xzxx10z1zzxz111000xxz001x0xxzxxzzxxzxxzxzxzzxxxxxzxzxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
