class c_184_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_184_6;
    c_184_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zxz00z0010zxx11zx00zxxz1zz100zzxzxzxzxzzxxzxzzzxxzxxxxzzxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
