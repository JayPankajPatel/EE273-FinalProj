class c_243_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_243_6;
    c_243_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0zzz01110x00xxx0x0x1xxzz0xxz1xzzzzxzxzzxxzxxzzxxzxxxxxxzxxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
