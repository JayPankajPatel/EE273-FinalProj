class c_82_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_82_6;
    c_82_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "001z0z0x100100z1111100xz1xx11101zzzzxxzxxxxxxxxzzxzzzxxzxxzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
