class c_881_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_881_6;
    c_881_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzx00x0z0xzx0xxz10xz1100xzxz11xxzzzzxzxxzzzzzxzxzzxxxzzxzzxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
