class c_1434_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1434_6;
    c_1434_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx1101xz0z00x01zxzxz1x0xzz0zx110xzzxxzxzzxzxzxzxxxxzxzzxzzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
