class c_1564_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1564_6;
    c_1564_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz00x0x1zx0zzz10100010001zzz10z1xxxzxxxzzxzzzzzzxxzxzzxxzzxzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
