class c_1039_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1039_6;
    c_1039_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0010z0zx10xz1xxx1x11110zzz01z0z0zzzxxzxzzzzxxxzzxxzxxxxzzzzxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
