class c_1664_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1664_6;
    c_1664_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx01z110x01x000xzxx0x100x10xx110zxzzzxzzzzxzxxzzzxzzzzxxxxxzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
