class c_1578_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1578_6;
    c_1578_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xxxxz1x10x11zzzx1zx010x11xzzz11xxzzxxxzzzxxzxxzzzzzxzzzzzzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
