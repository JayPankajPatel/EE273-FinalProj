class c_931_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_931_6;
    c_931_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x010z1z1zz1x00x0zxx10x10zz011z0xxzzzzxxxzxzxxzzxxzzzxxxxxxxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
