class c_1318_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1318_6;
    c_1318_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0zzzzxz01xz1xx11z0zz11x0011xxx1zzxzzzzzzxxzzxxxzzzzzxzxzxzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
