class c_1316_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1316_6;
    c_1316_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z111xzz01x1001zzzz1011xz00z0zxxxxzxzzxzzzxxzzxzzzxzxxxxxxxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
