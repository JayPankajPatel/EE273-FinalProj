class c_1667_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1667_6;
    c_1667_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1zxzx1xx10z0x0zzxz001zx00z1xxx0zzzxxxzzzxxxxzxxxzzxzxzxxzzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
