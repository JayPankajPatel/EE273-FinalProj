class c_1488_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1488_6;
    c_1488_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z0x1xzz0xz110zzz0zzxxxz1z01z011zxxxzzxxxzxzzxzzxxzxzxzzzzzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
