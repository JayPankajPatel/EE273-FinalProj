class c_438_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_438_6;
    c_438_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x01xxzzx1zzx1z1z01x1011zz01x110zzzzxxzzxxxzzzzxxxzzzxxxzzzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
