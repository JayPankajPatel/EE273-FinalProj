class c_1245_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1245_6;
    c_1245_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "100z010x01zx1xzz10z0xxz1z001x0x1xxzzxzxxzzzxzzxzzxxxxzzxzxzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
