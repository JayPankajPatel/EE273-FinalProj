class c_887_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_887_6;
    c_887_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zxxxx0110x001xz0xxzx11x0z00x01zxzzzxxxzxzzxxxzxzxxxzxzxxxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
