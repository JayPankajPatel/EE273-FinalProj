class c_1705_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1705_6;
    c_1705_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11xxxzz10x1zzzxzzzz1x0x100xz1z10xxxzzxzxzzzzxzzxzxzxxzxzzxxxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
