class c_631_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_631_6;
    c_631_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxz0zx10xzxxzx1zzzxxzz0z01x10zx0xxzxzxzzzzxzzzzxxxxzzxxzzxzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
