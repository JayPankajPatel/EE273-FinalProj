class c_1293_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1293_6;
    c_1293_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zz1z11xxx0zx0zx0xxx0zzx01z0z00xxxxzzxxxzxzxzxxzxzxzxzxxxzzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
