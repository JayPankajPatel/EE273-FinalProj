class c_1530_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1530_6;
    c_1530_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z00001011x10x0x11x00z0x1z0xxz1xzzxzzxzxzxzxxxxzzzxxxzzxxxzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
