class c_48_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_48_6;
    c_48_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11x1xzx0z0xxxzzx110001zz0000111zzzzzxzzxxxzxxxzxxzzxzxxzzzxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
