class c_707_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_707_6;
    c_707_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1101xxzz0xzzx1xz1x1xxz01xzz1111xxxzzxzxxxzxzzxxzxxxzxzxzxzzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
