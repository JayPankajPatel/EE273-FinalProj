class c_596_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_596_6;
    c_596_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01xx0z0xx0x101z10z00000xx011z0zxxxxxxxzxzzxzxxzzzxxzzzxxxzzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
