class c_1741_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1741_6;
    c_1741_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1011z01z01010z00xxzx1z11xx010001xzxzzzzxxzzzxzxzxxxzxxzxxzxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
