class c_873_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_873_6;
    c_873_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1xz11z0z011xxx1zzzz10z110z0xxx1xxzxxzxzxxxzzxxzzzzxxzxzzzxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
