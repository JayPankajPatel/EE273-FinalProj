class c_1498_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1498_6;
    c_1498_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0zzx1zxx100xx1z0x0xx0x11xz10z10zzzxxzxzxxxxxzzzzzzxzxzzzzxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
