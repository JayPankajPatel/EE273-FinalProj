class c_811_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_811_6;
    c_811_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01x0z00000z01zzx10x11zz1100zzxx0zzxzzxzzzzzzxxzxxzzzzxxzxzxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
