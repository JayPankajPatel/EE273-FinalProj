class c_1170_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1170_6;
    c_1170_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1z1xxx0zz0xxxzzz0xz1z0zx0z10x11zxxzxxxzzzxzzzxxzzzzzzzxzzzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
