class c_679_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_679_6;
    c_679_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0zz1z10xzx0xzx10x01z0z110zz000xxxzxxxxxzzzzxxxxzzxxzzzzxzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
