class c_603_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_603_6;
    c_603_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0z00xz0111z100x10zzx11xzx010z10zzzxxxzxxzzxxzxzzxxzxzzzxxxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
