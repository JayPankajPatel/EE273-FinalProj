class c_846_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_846_6;
    c_846_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x1010zzzzz101011z1zz1001zxz1zxxxxzxxxxzzxxzzxzzzxxzxzxxxzzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
