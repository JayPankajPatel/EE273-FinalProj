class c_938_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_938_6;
    c_938_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z01xzzxx111111zzz00010zxx0xzz1x1zzxxzzzzzzzzzxzzzxxxzzxxzzxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
