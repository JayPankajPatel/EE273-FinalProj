class c_929_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_929_6;
    c_929_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z11x00z1xx1xxxxxxx010zz0xzz0zxxxxzzzzzzxzzxzzzzxxzxxzxzzxzxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
