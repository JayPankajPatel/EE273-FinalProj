class c_56_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_56_6;
    c_56_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z1z0xz100x1xxzxx1zxzzx0010z1zxxzzxxzxxxxzzzzzxzzxzzxzxxxzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
