class c_1506_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1506_6;
    c_1506_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzz0x0z0xxxx00xz01z0zz11x0z00zz0zzxzzzxxxxxzzzxzxzzzxxxzzxzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
