class c_861_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_861_6;
    c_861_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11zx100x0111zxz1x0x1x10z1x00010xzxzxzzzzzxxxzzxzzxxxzzxxzzzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
