class c_1095_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1095_6;
    c_1095_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "110zzz0x0101z00xz00x111010111011xzxzzzxzzzxzzzzzxxxzxzzzxxxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
