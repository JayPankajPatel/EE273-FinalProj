class c_1341_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1341_6;
    c_1341_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx1xx1zz1xz1101z00001zzz11x00zxxxzxxzxzxzxzzzzxxzzxzxzzxxzxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
