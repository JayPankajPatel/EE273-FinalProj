class c_1047_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1047_6;
    c_1047_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11z0xz0xx1zx010zx10101z10z0z1x01xzxzzzxxxxxxzzxxxxzxzxzzzzzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
