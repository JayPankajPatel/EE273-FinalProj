class c_1768_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1768_6;
    c_1768_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zzxx01x0xzxx0x0zx1x0100x00zzz01xxzzzxxzzzzxxzzxxzxzxzzxzzxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
