class c_1812_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1812_6;
    c_1812_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z1x11xx01z11x1xz1000zx01zx1z101zxzxxzzxzzxzzxxxzzxxzxzzxzzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
