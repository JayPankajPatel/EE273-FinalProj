class c_1296_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1296_6;
    c_1296_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0000x0x1zz01zx110x00z10xx10xxzzxzzxzzzxxxxzzzzxzzzzxzxzxzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
