class c_277_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_277_6;
    c_277_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1101zzxx11xx10z010110xx00x000101xxxxxzxzxxxzxxzxzzzzzzzzxxxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
