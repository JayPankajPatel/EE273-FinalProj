class c_1128_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1128_6;
    c_1128_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111011zxz1zzxx11x0x110z1z101z1z0xxxzxzzzxxxzzzzzzzzzxzxzxxxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
