class c_716_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_716_6;
    c_716_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zx000z110z1zz11x01zxx1z100x0zz0xxxxxxzzzxxzxxzxzzzzxzxzxzzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
