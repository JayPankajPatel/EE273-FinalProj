class c_1660_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1660_6;
    c_1660_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1x1x00xx00xz1zz0x1zxz0x0x1z001xxzxxzxxzxzzzxzxxxxzzzxxxzxzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
