class c_866_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_866_6;
    c_866_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "101x1z00xxz01xzz0z01xzz11zzxxzzzzxxxxxzxzxxzxxzzzxzxzzxxzzxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
