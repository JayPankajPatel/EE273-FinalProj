class c_1251_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1251_6;
    c_1251_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx0zz0x11100z01zx00z1100z1zz11z1zxzzzxxzxxxzxxzzxxzzzzzzzxxzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
