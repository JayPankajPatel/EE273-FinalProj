class c_961_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_961_6;
    c_961_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzx01z01x0z11010zxz00zxx1z10xx1zxxxzzzzxxzzzxxzxzzxxxzzzzzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
