class c_469_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_469_6;
    c_469_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z00x11z011z110x1x111zx0x0x1x1110xxzxzxxxxxxzzzxzzxzxxxzzxxzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
