class c_1865_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1865_6;
    c_1865_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1000x1x0x11z1xzxz00xzzz0001zxxzxzzxzxzxxzzzxzxzzxzzzzzxzzxzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
