class c_937_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_937_6;
    c_937_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1110x0z001x111xzzz0101xxxx00z1xzxzzzzxxzzxxzxzzzxxxxxzzzxxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
