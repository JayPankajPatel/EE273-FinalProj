class c_853_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_853_6;
    c_853_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zz1xxz00z001x1z0011xzzz10zz1zz0xzzxzxxxxxzzzxxxxxxzxxxzzzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
