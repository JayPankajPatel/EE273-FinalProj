class c_176_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_176_6;
    c_176_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xzz1zz1110z0011zxxxzz11zxx0z00zzzxzxzxzzzxzxxxxxzxxxzxxzzzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
