class c_800_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_800_6;
    c_800_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01xzzx00x00xz111x00xxzz0x01x0z00zzzzxzzxzzxxxzzzxxxzxzxzzzzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
