class c_1417_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1417_6;
    c_1417_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0111z0x0zxz1011zxx0xxzxx111xxzzzxxxxzzxzzxzzxzzxzzzxzzxxxxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
