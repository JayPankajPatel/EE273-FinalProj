class c_1068_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1068_6;
    c_1068_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1xzxx1x1xz1x101zz11111x1zx1xzz1zzzzxxzzxzxxxzxxzzzzxxxxzxzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
