class c_1465_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1465_6;
    c_1465_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "000z0x0xzx1z00z0z01zzx011x011011xxxzzzxxxxzzxzxxzzzzxzzzxxxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
