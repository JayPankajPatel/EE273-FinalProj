class c_1201_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1201_6;
    c_1201_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xxzzzz101zz10x110xxzz1x0z0zxx11xxzxzxxxxzxxzxzzzzxzxzxzxxxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
