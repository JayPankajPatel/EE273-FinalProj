class c_1873_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1873_6;
    c_1873_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx111xx10z0x1xxzzxz111xz01zz01x1xxxxzzzzxxxxxzzzxxzxzxzxxxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
