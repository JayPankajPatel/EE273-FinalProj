class c_1677_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1677_6;
    c_1677_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1xzz11zx11zx100xxzxz1zzx1x0zzx0zzxxzxzzzzxxzxxxzxzzxxxzzzzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
