class c_1115_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1115_6;
    c_1115_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z01xx10xzz10x0x1xx00xxzz1z0z001zzzzzzxxzxzzxzzxxxxzzxxxzzxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
