class c_1491_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1491_6;
    c_1491_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzxz0z1010x01z100xx10zxz10zz00xzxzxxzzxzxxxzxxxxxzxxxxzzzxzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
