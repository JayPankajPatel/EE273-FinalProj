class c_1694_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1694_6;
    c_1694_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x101x10xx0z111xx0zzz0110xx1z0001xzxzxzzzzzzxxzzzzzzzxzzzxzzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
