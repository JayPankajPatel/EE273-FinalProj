class c_34_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_34_6;
    c_34_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1z1001011x1xx11xxz0xx0z01z11x10zxzxxxzzxxxzzxzxzxxzzzzzzzxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
