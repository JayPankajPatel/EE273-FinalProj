class c_1136_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1136_6;
    c_1136_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1xzz0x0zx0x1x00z10x0xxxxx1zz0xzxzxzxxxxzzxzxzxzzxzzzxxzxxzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
