class c_902_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_902_6;
    c_902_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zzzx11xx10010111xx110zzx0x111xxxxxzzxzzzxzxzzxxzzzxzzxxxxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
