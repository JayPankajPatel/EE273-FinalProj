class c_109_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_109_6;
    c_109_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzzzxzx110x01xxxz01zz100xxx1xx11xzxzxxzxzzzzxxzxzxzzzxxzxzxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
