class c_1584_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1584_6;
    c_1584_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x01xxx1000x0z01z10x01zx0z0zx1000zxzxzxzxzzzzzzzxxzxzzxxzzzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
