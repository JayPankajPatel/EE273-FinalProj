class c_1566_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1566_6;
    c_1566_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx00xz0z01x0zz10zz10xz0100xzz000xzxzzxzzzzxzxxxzxxzxxxxxzxzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
