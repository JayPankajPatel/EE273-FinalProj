class c_1072_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1072_6;
    c_1072_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z10zz010xzx00zz0x110x0xxzxx0xzzxzxxzxxxzxxxzzzzxzzzzxzzxxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
