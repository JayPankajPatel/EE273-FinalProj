class c_1558_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1558_6;
    c_1558_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z11zxzxx1xzzz00001x0z0xz1z1z0010zzzzxxzxzxzzxxzxxzxxxzxxxxzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
