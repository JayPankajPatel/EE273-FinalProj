class c_443_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_443_6;
    c_443_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz000xzx1xzx1z001z0xz10zx0zx10x1xzxzzzzxzxzxzxxzxzxzxxxzzxxzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
