class c_535_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_535_6;
    c_535_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1zxz100x1z1z11zzz0xzz1x0z0z110zzzxxzzxzxxxxxzzzzzxzxxzxxxxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
