class c_1458_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1458_6;
    c_1458_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzxz00zz1x11x11xx00zz0zxxx1zz11xxzxzxxzxxzzzzzxxxzzzzzxxxzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
