`ifndef __TB_PKG
`define __TB_PKG
`include "uvm_macros.svh"
package test_pkg; 
    import uvm_pkg::*; 
    // put includes here
    `include "tb_agent.svh"
    `include "tb_env.svh"
    `include "tb_test.svh"

endpackage : test_pkg
`endif // __TB_PKG 
