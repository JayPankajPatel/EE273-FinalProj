class c_1130_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1130_6;
    c_1130_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxxzz0zzxzxxz0z1zz0001z1z101xx01zxzxxxzzzxzzzxzxxzzxzzzzxxxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
