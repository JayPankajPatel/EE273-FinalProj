class c_1634_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1634_6;
    c_1634_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "110x0zx0x10z00xz0z0x00zxx0zz1x0zxzxzxzxxxzxxxzzzxzxzxzzzxzxzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
