class c_1617_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1617_6;
    c_1617_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx01x1z010zz001x0z01zx0zz0x10zxxxxzzzzxxxxxxxxzxxxxxxxzxzzzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
