class c_1523_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1523_6;
    c_1523_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzz11xzz11zx0z1zz10z10xz01zx00xxxxxxxxxxzxxzxzxzzzzzzxzxzxxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
