class c_1615_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1615_6;
    c_1615_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1z1xz0z0zzzx1xzx0xzzx1xxzx0zzzzzzxxzzzzxzzxxzzzxzxzxxxxxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
