class c_859_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_859_6;
    c_859_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00101z1xxx00zzzzxz101z10z1111101xzzxzzzzxxxzxxxzzzxxxxxzzxzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
