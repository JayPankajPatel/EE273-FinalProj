class c_854_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_854_6;
    c_854_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz1z01xz1xx10xzxxzz10z11101x11z1zxxzxzzzzzzzzxxxzzxzxzzxzxxzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
