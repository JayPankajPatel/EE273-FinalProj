class c_597_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_597_6;
    c_597_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0xx0zxzzzx110x111zz101xxx1zx1xzzxxxxxzxxzzxzzzzxzzzzxzzxzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
