class c_454_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_454_6;
    c_454_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1xxxx11101xx00x1010011z101z101zxxzxxzxxxzzzzxxxzxxxxzxzzzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
