class c_1446_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1446_6;
    c_1446_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10xxz10xxxx0z0zxx100zx10001xxxzzzzzxzxzzzxxzzxxzxxzzxxxzxzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
