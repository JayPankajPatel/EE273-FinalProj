class c_1621_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1621_6;
    c_1621_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0z10z11xz111xzxzzz01xx0xz110x11xzxzxzxzxzxzxxxxxxxzxzzxzxzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
