class c_959_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_959_6;
    c_959_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1110zzxz0z1x01xx00zzxz0111z101xzzxxzzzzxxzxzzxxzzxxzzzzzzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
