class c_676_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_676_6;
    c_676_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xz000111xz1xz01zz0xxxxx0xzx0xx0xxxxzzzzzxzzxzxzxzzzxxxxxzzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
