class c_700_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_700_6;
    c_700_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01110z1100x110zz01xz0z11zzzzzxxxzzxxxxzzxzzzxzxzzxxxxzzzxzzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
