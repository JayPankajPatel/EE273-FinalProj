class c_1724_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1724_6;
    c_1724_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z11zxz0x100z0zz0xxx0011zzzz00x1zxxxxxzxzxxxxxzxxzzzxzxxxzzzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
