class c_144_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_144_6;
    c_144_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0111z00x1xxz1xzzz00x1011xxz11100zxxzxxxxzxzxzxzzxxzzzxxxxxzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
