class c_1783_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1783_6;
    c_1783_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzxxx111z1zzzzx0zx001z101zz0xz10zzxxxxxzzzzxzzzzxzzxxzxxxxxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
