class c_437_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_437_6;
    c_437_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z010x111z0zxz00001z00z1z1101xzzxxxzzzxzxxzzxxxzxxzxzzxxzxxxzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
