class c_727_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_727_6;
    c_727_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00zzx00xxz11xz11x00z0x00xzz0000zxxxzxxxzzzxzzzzxxzzzxzzzzzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
