class c_549_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_549_6;
    c_549_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0xxz1zzxz10xz1z0x1x0xxz0xzz001xxzzxzxzzxzzxzxxxzxxzxzxxxzzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
