class c_1228_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1228_6;
    c_1228_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0zxx0z1z01x1101xx001xx001z0zzz1zzxxxzzxxzzzxxzxzzxzxzzxxzxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
