class c_214_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_214_6;
    c_214_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zxx11x1zxx1x1z1z0z11x0x1zzx0zz1xxzxxxxxzzxxxxxxxxxzxzzxxxxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
