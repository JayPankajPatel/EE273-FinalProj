class c_1652_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1652_6;
    c_1652_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1z1zz11zz0x0101xzzz1x1xz10xz1xxzzzzxzzzxzzzxzzxxxxzzxxxxxzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
