class c_684_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_684_6;
    c_684_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xzzxzzzz00z000z00x00x0z00zz1xz1xxzxzxzzzxxxzzxxxzzzxxxzzzzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
