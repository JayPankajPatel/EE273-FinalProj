class c_1593_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1593_6;
    c_1593_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1xxzzx001z0z1zxzxxz0010x01x100zxzzxzxzzzxzxzxzxzxzzzxxzxzxzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
