class c_1057_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1057_6;
    c_1057_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzxxz1xxz0zxzxz111x0zxzzxz111xz0zzxxxxzxxzxxzxxzxxzxzxxzzzzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
