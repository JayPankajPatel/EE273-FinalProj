class c_726_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_726_6;
    c_726_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "001xzx10000z0zxzz1101z0xx10z1z1zxxxzzxxxxxzxxzzzxzzzxzxxxxxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
