class c_864_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_864_6;
    c_864_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10zxxx0z0zx000xx001001xxxzxz1x0zzxzzzzxzzzzzzzzxxxzzzxzxxzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
