class c_1730_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1730_6;
    c_1730_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz1x0010zz1zzxz0001xz1xz0x001zxzxzxzzzxzxxzzxzzxxzxzxzxxxzzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
