class c_463_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_463_6;
    c_463_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0z11z01z101z1x100z11x110zzxz0xxzxzzzxxzzxzzxxxzxzzxzxxxzxzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
