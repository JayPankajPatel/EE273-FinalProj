class c_614_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_614_6;
    c_614_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0xxzz001x01zxxxz001000xz001zzzxzxzxzzxxxxzzxzzxxzxzzzxxxzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
