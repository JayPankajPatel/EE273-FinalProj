class c_1131_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1131_6;
    c_1131_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx1x101110x0x0xx1xx001x011x0zz1xzzzzxzzxxzzxxxxzzxzxzzxzxzzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
