class c_1363_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1363_6;
    c_1363_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0xxx101zzz101zz1z0z101xzxxx010xxxzzxzzxxzzzzzzxxxzzxzzxzxxzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
