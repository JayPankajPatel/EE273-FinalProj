class c_282_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_282_6;
    c_282_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzxxz10z01z0x01x1xxzz1111zxx11zzxxxxxzzxxzxxzxxzxzzxxxxzzxzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
