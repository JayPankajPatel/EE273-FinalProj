class c_441_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_441_6;
    c_441_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0xxxzz1zxxx1z10110z11010x0x100zzxxzxxzzxxxzxxzzxxxxzzxzxzxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
