class c_1736_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1736_6;
    c_1736_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx0xzx1zxxx101zz0x1z1zz1x1z10xxxxzzxxzzxzzxzxxzxzzxzxzxxxzxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
