class c_1069_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1069_6;
    c_1069_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10zz01xz10zzx1xz1xxzxxx1xx10z1zzzzzzxxzxxxxxxxzzxxzxxxxxzzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
