class c_93_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_93_6;
    c_93_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10zxz01xz11zz1111xx1010x011zzxz1xzzxzxzxzxzzxxxzxzxzxzxzzzzzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
