class c_1688_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1688_6;
    c_1688_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zxx0zz010xx01z01x111z1zzxz1z00xxxxxxzzzxzxxzzxxzzxzzxxxzzxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
