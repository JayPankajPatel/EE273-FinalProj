class c_1258_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1258_6;
    c_1258_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx000z111x1z11100z1xx10x0z100zzzxxxzxzxxzxzzxzxxzxxxxzxxxzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
