class c_121_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_121_6;
    c_121_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z01zx11xz001zz10zxx1x01x01zzx0xxxxxzxxxzxxzzzzzzxxxzxzxxxxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
