class c_657_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_657_6;
    c_657_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz10z0011x0z1zxz11xz001z1z010zzzxxxxzzzzxzzzzxxzxzzzxzxxzzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
