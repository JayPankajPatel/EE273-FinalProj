class c_1771_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1771_6;
    c_1771_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x11x0z100zxxzx10xz0z1zx0zxx1zzzxzxzxzzxzxxxxxxxzxzzzzxzxzzzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
