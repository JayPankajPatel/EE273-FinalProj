class c_379_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_379_6;
    c_379_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z11zx1z000xzx00x111xx0z1x1x1xzzxzzzzxzxxzxzzzzzxzxzxxzzzxxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
