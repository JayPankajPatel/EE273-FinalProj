class c_780_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_780_6;
    c_780_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x0z11z10101x0101xzxzz01110x1xxxzxzzzzzxxzxxxxxzxxzzzzxzxxzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
