class c_1354_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1354_6;
    c_1354_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxxx0011x010x0x0zxx0xzxxxx00xx10zzzzzxxxxxzzxzzxxxzzzxzxzxzxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
