class c_741_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_741_6;
    c_741_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x10zxz1zxzz0111xzx1z10xxzzzzx1zxzxzzxxzzxxzxxzxzxxxzxxxzzxzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
