class c_650_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_650_6;
    c_650_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zzzxx0xz0x0x011zxxzx1x1100x0zx0zxxxxxzxzzzxxxzxxxzxxzzzzxxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
