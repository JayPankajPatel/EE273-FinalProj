class c_1281_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1281_6;
    c_1281_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0zx111xx01z1z10zzzz0xzx1z01xzx0xxzxzxzzxxxxxzzzxzzxzzxxzzxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
