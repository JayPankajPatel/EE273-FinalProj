class c_19_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_19_6;
    c_19_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1xz1100xx00zz11001x111z11xz101xzzxxzxzzzzxxzxzxzzxzzxxxzxzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
