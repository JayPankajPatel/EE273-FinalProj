class c_258_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_258_6;
    c_258_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x0z1z1zz0z0xx11xxx0z110x1zx0xxzzxxzzxxxxxxxxzxxxxzzxxzzzzxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
