class c_910_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_910_6;
    c_910_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1xz0z0zxzzxz1xx10zzzz10zzz01x11zzzzxzzzxzzxxzzxzxzxzxzzxzzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
