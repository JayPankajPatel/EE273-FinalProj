class c_1518_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1518_6;
    c_1518_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xzz10xz1x0xxx00xz1zx1xx100111xxxzxzxxxxxzzzxxzzxzzzzxzzxxzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
