class c_234_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_234_6;
    c_234_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zzx0zzz0011x1xxzz1zz001xz1101xxxzxxxzzzzxxzxzxzzxxzxxzxxxzxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
