class c_729_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_729_6;
    c_729_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z011z1z00zx10zzxx1z0zz1z0x0xx0z0xzzzzzxxzzxzxzzxzzzxzxzzxzzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
