class c_536_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_536_6;
    c_536_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11x111x1z1z0x01zzzz01000xz1zxzx0zxzzxzxxxzxzxzxzzxxxxxxzzxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
