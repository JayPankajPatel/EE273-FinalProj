class c_871_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_871_6;
    c_871_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxz0x1x10x101z110z1zx000xx110zx0xxxzxxzzxzzxxxxxxzxzzzxxzzxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
