class c_591_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_591_6;
    c_591_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z010xx0001x10z11xxxxxz011x011z0xxzxxxxzxzzzxxxxxzxxzxzxzzzzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
