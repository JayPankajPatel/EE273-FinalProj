class c_1089_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1089_6;
    c_1089_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x01z01zz0x0101xzzz00xxzx1z0zx0x1zzzzzxzxzzxzzzzzxzzzxzzzxzzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
