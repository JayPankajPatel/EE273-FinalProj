class c_1538_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1538_6;
    c_1538_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00x1z0010z000xzx0z0zzx1z00xx0x01xzxxzxxxzzzxzzzzxxxxxxzxzzxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
