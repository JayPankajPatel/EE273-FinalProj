class c_1426_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1426_6;
    c_1426_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1xzz1z0x1z1101z1z00000zzxx11z01xxxzxxxzxzzxzzzxxzzzxzzxzxzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
