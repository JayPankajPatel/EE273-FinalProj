class c_1457_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1457_6;
    c_1457_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x11xz01zz10xzzxz11zx1z1x0x110z0xzxzxxxzzzxxzxzxxxxxzxxzzxxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
