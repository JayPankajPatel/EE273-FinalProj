class c_1515_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1515_6;
    c_1515_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0z1zzz1000z0xxzz1xxx0zzz011zxx1xxxzxzxxxxzxxxxzxzxxzzxzzzzzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
