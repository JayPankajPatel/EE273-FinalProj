class c_28_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_28_6;
    c_28_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxxzxzxxx11zxzx0xx1xx10zx1xx10zxxzzxxxzxxxzzxxxzxzzzzzxxxzxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
