class c_1767_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1767_6;
    c_1767_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzz0x0zxz1x1zzxx111zx1z1z01z11zxxxzzxxzzxzxxxxzxxxzzxzxxzxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
