class c_956_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_956_6;
    c_956_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z00z0x0zxxxz00z00xz0xxxzxz100x0xxzxzxzxxxxzxzxxxxzxzzzxzzxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
