class c_228_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_228_6;
    c_228_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zz00z1x10xzz0x00zx0x0zzz10zzz0xzxxxzzxzzxxzxxzzzxxzxzxzxzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
