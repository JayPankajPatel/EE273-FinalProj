class c_658_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_658_6;
    c_658_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111xxx1010zxxxzz0x00z100xzxx1z0zzxxzzzxxzzzxzxzxxzzzxzxzzxzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
