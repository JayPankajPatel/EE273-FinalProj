class c_1508_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1508_6;
    c_1508_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z1x0xzz0zzz11xxzzz01z1x10z0z01zzxxxxxxzzzzzzzzzzxzzxxxxxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
