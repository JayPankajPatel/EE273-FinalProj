class c_989_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_989_6;
    c_989_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z01111xz00x10010zz11x0xz01z0xzxzxzxzxxzzzzxxzxxzxzxzxxxxzxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
