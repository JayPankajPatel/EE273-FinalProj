class c_1308_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1308_6;
    c_1308_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz10zz010x1xx10z0x01z1xx1111zx0zzxzzxxzzxzxxxzzzzzzxzzzzzxzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
