class c_1792_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1792_6;
    c_1792_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00z10xx01001011xx1zx0xxx001zzxz1xxzzxxxxzxzzxxxxzxxzzxxxzxzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
