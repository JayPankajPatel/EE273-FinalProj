class c_1053_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1053_6;
    c_1053_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z1z1xz1010xx1xx1zx0zx0xxx00x011xxzzzxzxzzxzxxzzxxxxxxxxxxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
