class c_265_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_265_6;
    c_265_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzx0z110zxz0z0010011zxx11zz11zz1zxzzzxxxzzzzzxxxxzzzzxzzzxxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
