class c_784_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_784_6;
    c_784_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10x10011x11xzz010xzz1xzz111xzxz1zxzzxzxxxzzxxxxzxxxxxzzxxxxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
