class c_1244_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1244_6;
    c_1244_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z10zx1x0x1zz0x0x1xx1101000x1zzxzzzzzxzzxzxxzxzzzzzzxxxxxzxxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
