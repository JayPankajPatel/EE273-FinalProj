class c_1352_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1352_6;
    c_1352_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11xxzz0z0010z1zxzxxx0z10000zxxx0xzzxzzxxzxxzzxzxzzzzzzxxzxxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
