class c_779_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_779_6;
    c_779_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1zz110xz00z0xzzz0x01zz0z0z1xxx1zzxzzxxxxxxxzxxzzzzxzzzxzzxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
