class c_1059_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1059_6;
    c_1059_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz110xxxxz0zz100zzz01x00z0zxz001zxxzxxxxzzzzxxxxzzzzxzzxxzxzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
