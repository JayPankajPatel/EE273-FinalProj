class c_1242_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1242_6;
    c_1242_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1x1z11zzz111x1x0x00000xx00x010xxxzzzzxxzxxxxzzxzzxzxzxzxxxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
