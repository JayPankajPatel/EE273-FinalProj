class c_1602_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1602_6;
    c_1602_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0x10x1x1x1101x0001zx1zz01100x11zxxzzxxzzzzzzxxxxzzzxxzzzxzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
