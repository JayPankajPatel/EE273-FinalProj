class c_1867_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1867_6;
    c_1867_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z001zzz0x001z011x0x01xxxzx0zx0z0xxxzzzxxxzxxzzzzzxzxxzzzzzzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
