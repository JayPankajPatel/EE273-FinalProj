class c_1322_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1322_6;
    c_1322_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzz11xx11z1zzxz1z0xz10x011000zz1xxzxxzzxxxxzxxxxxzxzxxxxxzzxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
