class c_791_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_791_6;
    c_791_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxx1x1zxx1100zx1000100x010x00zx1xxzxzxxxzxzzxxxzxxxxzzxxxzzzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
