class c_1713_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1713_6;
    c_1713_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zx1zx1z0x1x01zx01z1010x1x01z00zxxxzzxxzzxzxzzxzxzzzxxzxxxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
