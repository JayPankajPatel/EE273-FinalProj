class c_1217_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1217_6;
    c_1217_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10z1x0x1001101z0zxz1001x011xzxxzxzzxzzzzxzxxzxxzxzzxxxxxzzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
