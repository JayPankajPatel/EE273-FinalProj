class c_503_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_503_6;
    c_503_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0111xz0x1z11xzx1x01xxxz001x010zxxzxxxzzzxzzzzzxzxzxzzxzxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
