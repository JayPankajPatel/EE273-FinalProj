class c_92_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_92_6;
    c_92_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zxz01x1x01z11zzx1zz01z1z1xx1xz1zzzzzzzzxxzzzzxxxzxzzxxzxxxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
