class c_1794_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1794_6;
    c_1794_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zzzx0xxx1xx011zx0xz101z01z000zxzzxxzxxzxzxxxzxxxzzzxxxxzxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
