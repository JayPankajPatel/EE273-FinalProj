class c_771_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_771_6;
    c_771_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10x1zz1z111x0z0zx10x01z0zx01z0zxzxxxzxxxxxxzxzzxxxzxxzxxzzzxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
