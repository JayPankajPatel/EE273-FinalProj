class c_1527_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1527_6;
    c_1527_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00110xxzx00z0zz1x1xzx110z1zx1z0xxxzxzxxxzzzxzxzzzzzzzxxxzxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
