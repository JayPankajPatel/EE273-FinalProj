class c_313_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_313_6;
    c_313_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxz010xx0z0xzxxxzz010z1z00010xx0zzxxzxxxzxzzxzxzxxzzzzzzxzzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
