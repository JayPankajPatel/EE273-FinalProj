class c_295_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_295_6;
    c_295_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1xx0z0xz0x110z1xzx10zz0010z111zzxzzxzzxzzzzzzxxxxzzzxxxxxzxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
