class c_646_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_646_6;
    c_646_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "001x0xz1101xz01xx01xz0zzxzx10101zxxxzxxzzzxxzzxzxxzzxzxzzxxzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
