class c_816_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_816_6;
    c_816_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zx0x110zxz11xx101zx1x00xxx101zzzxxxzzxzxxxzzxxzxxxxzzzzzzxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
