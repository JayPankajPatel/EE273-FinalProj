class c_461_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_461_6;
    c_461_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0z0x0x1zz1xx11x1x0zxxz10xzzx0zxxzxzxxxzxxxzxzxzzxxxxzxzzxzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
