class c_1099_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1099_6;
    c_1099_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1110zxx1zx1x00zxzz0zx00zz00zxxxxzxzzxzzxzzzxxxxxzzzxzxxzxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
