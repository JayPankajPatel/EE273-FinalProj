class c_238_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_238_6;
    c_238_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10101x00xx0z11zz10zx001x110zzzxzxzzzzzxxzxzzxzxzzzzzzxxxxzzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
