class c_365_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_365_6;
    c_365_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x0xzz10xzxx0x0z101zxz0z1x0xzx1xzzxzzzzxxxxxxxxzzxzxxxzzxzzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
