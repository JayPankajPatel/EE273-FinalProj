class c_1196_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1196_6;
    c_1196_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "110000zzxx0z1z1zz101zx01xzxx1z1xzzzxzxzxzxzzzzzxxzxzxzxxzxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
