class c_1091_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1091_6;
    c_1091_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzx0111xx1zzz0zx011000111x0zz01zxxxxzzzzzzzzxxxzxxzzxxzxxxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
