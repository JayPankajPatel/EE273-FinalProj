class c_1863_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1863_6;
    c_1863_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0zz0z0z0z1z10zx01xz0z1xz10xz0xzzzzxxzxzxzxxxzxxzxzzzxxxxxxzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
