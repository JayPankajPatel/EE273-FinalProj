class c_1351_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1351_6;
    c_1351_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z11xxx1xz0z101xz1zxx10xz001x0001zzzxxxzzxxxzxzxxxzxzzxzzzzxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
