class c_1607_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1607_6;
    c_1607_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx1010x00z0z1xx00zzz00xxzxx0xz1xzxzxzzzxzxxxzxxxzzxzzxxxxzxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
