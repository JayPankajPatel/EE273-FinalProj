class c_998_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_998_6;
    c_998_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x0xx0x11z1z1zx11001xxzxxxx0x000zxxzxxzzzzxxzzzxxzxzzzzzzzzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
