class c_805_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_805_6;
    c_805_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxxxx10zxx1z11xx011001xz00110zz1xzzzzzxxxzzzzxzxxxzxxzzzzzxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
