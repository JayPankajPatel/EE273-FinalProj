class c_229_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_229_6;
    c_229_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10zxxxxxxzxzzz10x111zzz010x0x1zzzzzzzxzxzxzxzxxxzxxzxxxxzxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
