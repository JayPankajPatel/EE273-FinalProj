class c_129_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_129_6;
    c_129_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zz01011101xz0z1zx0001xxzx0x0zx0xzxxxzxxxxzxxzzzxxzxzxzxxxxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
