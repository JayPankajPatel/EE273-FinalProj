class c_668_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_668_6;
    c_668_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x0zz10zx0z11zxzzz11zz0110z0x101zzxzzzzxzzzzxxzxzzzxxxzzzxzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
