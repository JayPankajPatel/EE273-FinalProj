class c_756_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_756_6;
    c_756_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x11z11z0z0z01zzxzz01zzzzzzz1xxzxzzzzxzxzxxzxxzzzzzzzxxzxxxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
