class c_1204_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1204_6;
    c_1204_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1xz11xx11z0z10z1z11x0x1zz1x000zzzzzxxzxxxxzxxzzxzzzxxxzxxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
