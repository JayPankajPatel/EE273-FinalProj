class c_1490_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1490_6;
    c_1490_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x01x0z00x010zxz1zz1xx1z1000z1010xzxzxzzxxxzzxzxxxzzxxxzxzzxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
