class c_1103_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1103_6;
    c_1103_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzx1z00z0x01x0xxzxx1x10010x0zx11zzzxzzzzzxzxzxzxzzxxzxzzzxxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
