class c_396_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_396_6;
    c_396_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x100xz1zxx0zzxzxxz0x0zz001110z1zxxzxzxzxzzzxzxxxzxzzzzxzxxzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
