class c_863_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_863_6;
    c_863_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zzxz0x0z0z1xz111z01z0z000zzxz00zzzxxxxzxxzxxxxzzzxzzxzxzxzxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
