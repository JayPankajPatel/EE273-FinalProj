class c_528_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_528_6;
    c_528_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11z0zz011100xz1zxzxxzx100xz1011zxzzxxzxxxxzxzzxxxzxzxzxzzxzxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
