class c_1097_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1097_6;
    c_1097_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0xz110xz1z1xxx10z1z001xz1x1zxz0zzxxzxxzxzxzxxzxzxzxzzxxzxzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
