class c_1468_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1468_6;
    c_1468_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzxzx1011x0zx1zzx0zz0xx0x1x0xx11zzxxzzxxxxzxzxzzxxzxzzxxxxzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
