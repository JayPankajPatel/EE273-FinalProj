class c_1124_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1124_6;
    c_1124_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z11x1z0100xz0z0x1x0z0xz00x101z1xzzzxxzxxzxzxxzxxzzxzzxxzzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
