class c_1299_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1299_6;
    c_1299_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11zzx1xxx00zz0xxzxx001xzzxxx0z10xzxzzxxzzzzxxxzzxxzzzxxzxxxxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
