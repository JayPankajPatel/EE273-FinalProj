class c_1843_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1843_6;
    c_1843_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x0z01x0x1x1xzxzz1111zx0010001z0xxxxzxzzxzzzxxzzzxxxzzxzxzzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
