class c_1816_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1816_6;
    c_1816_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x1xxzx1110z10110z0z0xx1xx0101z1zzzxxzxzxzzzzxzxzzxxxxxxxzxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
