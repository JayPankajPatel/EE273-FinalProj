class c_1356_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1356_6;
    c_1356_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z10z10xx1x0xz101xz1z1xx1zx0x111xxzxxxxzxxxzxxzxzzzxzxzxzzxxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
