class c_1543_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1543_6;
    c_1543_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxx1xx0zxx10x1110x1z11xzxzx0zz11zzxxxxzzxxxzxxxxzzxxxzzzxxzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
