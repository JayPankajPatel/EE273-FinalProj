class c_696_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_696_6;
    c_696_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x1x0z1zxxx01z10x11001zx0xxxzz0xzxzzxxzxxxxxzzzxzxxzzzxzzxxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
