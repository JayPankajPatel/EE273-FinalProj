class c_1283_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1283_6;
    c_1283_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzx0xxxzxz0x110z101000111zx00xx0xxzzxxzzzxzxzxxxxzzxzxzxzzxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
