class c_384_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_384_6;
    c_384_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00x01xx10xxzzx01z0xz00z0xxz1x0zxxxxxzzzxzzzxxxzxzzzxxzxxzxzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
