class c_1166_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1166_6;
    c_1166_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0x1001z10z1z1zzzxz01x00010x000xzzzxxzxzzzxzxzzxzxzxxzzzxxzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
