class c_1532_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1532_6;
    c_1532_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10x1zxzxx100x0xx0011101z1zx1x1zzzxxzzzxzzxxzzzzzxxxzzxxzxxzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
