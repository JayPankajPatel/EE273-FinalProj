class c_1046_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1046_6;
    c_1046_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx1xzzxz1000xx10zx0xx00zzz0z11x0xxzzzzxzzxxxzzxzxxxxzzzzzxzzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
