class c_1671_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1671_6;
    c_1671_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11x0xzz0z001x11zx1z1z111z0xxxzz1zzxzxzxzzzzxzzxxzzxxxzzxzxxzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
