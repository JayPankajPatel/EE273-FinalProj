class c_1146_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1146_6;
    c_1146_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0z0zz01100zx0100111z00zzxxzz1zzzzxxzzxzxxzxzzzxzzzzxzzzzzzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
