class c_337_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_337_6;
    c_337_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10000z01xzx10x1x11011x10000xxzxxzxxzzzxzxzxzzxxxzzzzzzxzzzzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
