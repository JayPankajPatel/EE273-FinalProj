class c_917_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_917_6;
    c_917_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x00x10xzx0z10z110z0zz1z0z1z0zzzxzzxxzxzxxxxzzzxxzxxzxxzzxxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
