class c_1619_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1619_6;
    c_1619_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz1x00x1101zxzz0xxx1x110xxxxx100xxzzzzxxxzxzzxxxxzzxzzzxxzzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
