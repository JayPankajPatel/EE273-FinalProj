class c_1202_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1202_6;
    c_1202_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx100xzz1x0zzxzzzzxx0z1x10zz01x0xxxxzzxxxzzxzxzxxzzzzxxzxxzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
