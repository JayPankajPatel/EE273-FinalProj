class c_1290_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1290_6;
    c_1290_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz1zz1xx10zx0x101zxx1zz0xzx00xxzzxzxzzzzxxzzzzxzxzxzxxxzxzzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
