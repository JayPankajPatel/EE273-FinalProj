class c_212_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_212_6;
    c_212_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z1101zz00xzx1z101z11zx1z00x0zzxzxzxzzzzzzzxxxzxxzxzxzxzxzxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
