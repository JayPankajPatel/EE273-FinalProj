class c_418_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_418_6;
    c_418_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzz01z001z00zx0z01x001z11z0xx01xxxzzxzzxzzxxzzzxzxxxxzxxxxzzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
