class c_403_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_403_6;
    c_403_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zz11xz1001zz0z101x110xzzx0100xxxzxzxxxzzzzxxzxxzxzzzxxxzxzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
