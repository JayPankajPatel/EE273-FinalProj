class c_760_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_760_6;
    c_760_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "110z110xxzzz11zxzzx0z100z0zzxxzxxxxzxxxxxxzzxzxzxzxxxzzxzxxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
