class c_1743_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1743_6;
    c_1743_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00z00000xxxxz0zx10zz1xxz0x1zxxz1xzzzxxzzxzxxzxxzzzzxxzxzzzzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
