class c_817_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_817_6;
    c_817_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx1z001z10z110xxz0z0111zxxxxx001xxzxzzxzzxxzxzxzzzzzxzzzxxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
