class c_366_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_366_6;
    c_366_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz0x11zzzx01z11zxx1zx1x11000zz0xzxzzzxxxxxxxxzzxxxxxzxzxxxzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
