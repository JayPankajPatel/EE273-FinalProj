class c_1153_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1153_6;
    c_1153_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z00xz01zxx1x0zxzzx10z11101001z0zzzzzxzzxzzzxxxxxxxxxzzxzzxxzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
