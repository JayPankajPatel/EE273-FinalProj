class c_361_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_361_6;
    c_361_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzz1z110z01z1xz0xzzx0xxxzzxx01xxzzxxzxxxzxxxxzzzzxzxzxzzzxxzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
