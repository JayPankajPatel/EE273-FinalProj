class c_675_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_675_6;
    c_675_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzxz10zz1z0xxz11x00z01zz0000zz10zzzxxzxzzxxzxxzxxxzzxxxxzzzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
