class c_1624_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1624_6;
    c_1624_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z00x10zz010xxxzxxzzx0z1001xx1110zzzzzxzzxxzzxxzzzxxzxxxxxzzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
