class c_351_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_351_6;
    c_351_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01z1z010zx1x00zx01zx0zx11zxzzzz1zzzxxxzxzzzzxxzzzzxzzxzxxzzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
