class c_1856_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1856_6;
    c_1856_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10zz0xz0xz1x0zx0xz0xxxxxzzxzxxz1zxzzxzzxzzxxzxzzxzxzzzxxxxzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
