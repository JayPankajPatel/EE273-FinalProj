class c_975_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_975_6;
    c_975_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x010x1z0xz11x00xzzz11x1xxz011z0xxxzzzzzxxxxzxxxxxxxxzzzxzxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
