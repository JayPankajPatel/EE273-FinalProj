class c_1851_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1851_6;
    c_1851_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0x00z0100xxx11x0x11xz100zxxx1zxzxxzzxxxzzxzzxzxxzzxxzxzxxzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
