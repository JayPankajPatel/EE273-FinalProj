class c_1052_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1052_6;
    c_1052_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzzx01xxx11z1x10zxz00zzxz000xz00xxxzzxzxxzxzxzxzxzxxzxxxzxxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
