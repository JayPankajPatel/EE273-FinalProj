class c_64_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_64_6;
    c_64_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10x0x0xzz00z0z01zzxzxx111z1zxxxzxxxxzxxzxxzxzzzzxxzzzxzzzzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
