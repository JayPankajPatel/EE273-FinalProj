class c_133_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_133_6;
    c_133_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0zxzxxzzx110zzx0111z1x110xxz1xxzxzxxxzzzxxxxzzxxxxxxxxzzzxxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
