class c_1839_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1839_6;
    c_1839_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10zzx0x00zx1xzz001z0xxz111zz0z0xzzxzzxxzzxxxzxxzzzzzxzzzzzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
