class c_1579_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1579_6;
    c_1579_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01z0001x1000010z1x110z1z0100x1zxzxzxzxzzzxzxzzxzxzzxxzxzzzxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
