class c_180_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_180_6;
    c_180_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1010z1xx1zxz010zz1xz01xz01010000zzxzzzzxxxzzzxzxxzzzxxzzxxxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
