class c_6_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_6_6;
    c_6_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "010z010zzx0x00z10zxx0zz100x0z0z0zzzzxzzxzzzxzzxzxxxzxxxzzzzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
