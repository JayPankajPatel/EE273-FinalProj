class c_1651_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1651_6;
    c_1651_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zxzx00x1xxxz0101z1111xzz0z010xzzzxzxxzzzzzzxzzxzzzzxxzzxzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
