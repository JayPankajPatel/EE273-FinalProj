class c_1706_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1706_6;
    c_1706_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzx00xxx11x10zz100z1xz1z0x00zz10xzzxxxzxzzxxzzzxzxxxzxzxzxzzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
