class c_1291_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1291_6;
    c_1291_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1011xzx00xzz1x0zzx10xzxzzzxz1x1zxxzxzxxzzxzxxxxzzxzzxxzzzzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
