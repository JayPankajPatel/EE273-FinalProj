class c_45_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_45_6;
    c_45_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1zxx110x1x1zzz101zz010xxz1zx0zzxxzxxxxzxzzxzzzzzxzzxzxzxxzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
