class c_1613_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1613_6;
    c_1613_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "000zx111xzzx100z00x1x0z1110xxzxxxzzxzxzzxxzzxxzzxzzxxxxzxzzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
