class c_1173_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1173_6;
    c_1173_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxxz0xx100xzxzx000xx0x1z1z01zx00xzzzzzzxzzxxxxxzxzxxzzxxzxxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
