class c_77_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_77_6;
    c_77_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11xzxxzz0xz1x001xzz101z0xz1zxzx1zzxxzxzxxxzzzzxxzzxxzzxzzxzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
