class c_1150_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1150_6;
    c_1150_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0xx1z0xz01z0x01zz00z0x10zzxz0zzzzxxzxxxxzxxzzzxxxzzxxxzzxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
