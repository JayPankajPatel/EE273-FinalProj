class c_294_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_294_6;
    c_294_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0z000001z01zzz00z0zx0xz100z100xzzxzzxzxzxzxzzzzxxzxzzzzzzxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
