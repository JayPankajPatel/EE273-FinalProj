class c_831_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_831_6;
    c_831_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "011zzxxxxx10x00xx1zz110x10zzzxxzzzxxzxzzxxzxxxzxzxzxxzzzzxzxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
