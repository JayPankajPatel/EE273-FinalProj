class c_301_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_301_6;
    c_301_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz1x111xzx0zz0x10z0x00zxzx0xz001xxzxzzzxxzxxzxxxxzxzxxxxxxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
