class c_1269_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1269_6;
    c_1269_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x11xx0xz00110z01zx0xzxz01z1z101zzzzzxxzzzxxxxzxzzxxxxxzzxzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
