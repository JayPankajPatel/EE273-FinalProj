class c_1029_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1029_6;
    c_1029_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzzxz111xxz0000z0xxzx1x1zx001zz0zxzzxzxxzxzzxzzzxzzzzxzxzzxzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
