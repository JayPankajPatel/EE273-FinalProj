class c_1763_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1763_6;
    c_1763_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111zx01xxxxx0zzx010001x0z1x10000xxzxxxzzzxzxxxxzxzxxxzxzzxxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
