

function tr_msg sb_predictor::sb_calc_exp(tr_msg t);
    // not implemented yet
    `uvm_info("Ref Model", "not implemented", UVM_LOW)
endfunction : sb_calc_exp
