class c_363_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_363_6;
    c_363_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0zzx1zxx11xz1x1zz01x1xzx0001z01xzzxzzzzzxzzzzxxzxzxxzzxzxzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
