class c_1701_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1701_6;
    c_1701_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x0x0z10zzx0010z0xz110zz0110x000xzxzxxzzzxxzxxxxzzxxxzzxxzxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
