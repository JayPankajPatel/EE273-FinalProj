class c_24_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_24_6;
    c_24_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xzx0x1111zzxx101xz1x100z000x10zzzzzxzxzzzxzzzzzzzxzzxzzxxzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
