class c_778_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_778_6;
    c_778_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x01x0z1xxzx1xxx1x11zzz1xz1x10x0xzzzxxxzzzzxxxxxzxxxzzxxzzxzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
