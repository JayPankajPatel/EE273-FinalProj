class c_1048_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1048_6;
    c_1048_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "000xx1110x1011zxxz0xzzx1zzx00101xxzzzxxzzxzzzzxzxxzzxxzxzxzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
