class c_935_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_935_6;
    c_935_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzxx110x010x010zz01xz010x1z1zz01zxzxzxzzzzzzxxzxxxxzzxzzxzxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
