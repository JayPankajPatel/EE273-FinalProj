class c_134_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_134_6;
    c_134_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz00zzzz1xxzzzz0xx0z10xz1z010zxzzzxxxzxzxzxxxzzxxzxzzxzzzzzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
