class c_412_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_412_6;
    c_412_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zxz0x1xzz01z0x0zx1zzzx1zxzz0zxxxzxxzzxzzzzxxzxxzzzxzxzxzxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
