class c_1815_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1815_6;
    c_1815_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0x00x01x1xx111z00zx1zx0zzzxx0zxxzxxxzxzzxxzzzzxzzzzxzxzxzxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
