class c_286_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_286_6;
    c_286_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz00z1x0z0x11x0xzx011z0xz10z00z0zxxzxzzzzzxzzxxzzxxzxxzzzzzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
