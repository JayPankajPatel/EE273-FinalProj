class c_1278_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1278_6;
    c_1278_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxz11010z01z0z10z100xx000100xx00xzzxzxzxzxxxzzzzxzzzzxzzzxzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
