class c_1385_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1385_6;
    c_1385_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00x11001x0x0111x011z1x0xxzzzzzx1xzzxzzzzxzxzxxzzzxxxzxxxxxxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
