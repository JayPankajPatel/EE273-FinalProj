class c_1809_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1809_6;
    c_1809_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzxzx1z00101101z1zx0z00zz1z01zx1zzxzxzzxzxxzzzzzxzxzzxxzxzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
