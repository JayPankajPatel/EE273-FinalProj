class c_615_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_615_6;
    c_615_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1001101x0x0101z0xxz11100z0zx1z1zxzxxzxxzxzzzzzzxxxzzxxzxzzzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
