class c_1197_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1197_6;
    c_1197_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xx1xz0zz1z000xzx01x0z00xz0z1xx0xzxzxxxxxxxxzxxxzxxxxxzxxzzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
