class c_1514_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1514_6;
    c_1514_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x001111z1xzx01xx100zzxxz0z0zx0z0xzxzzzzzxxzxxxxzxxxxxxzxxxzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
