class c_1234_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1234_6;
    c_1234_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxx1xz1xx10x1z110xxxz0010x110zz1zzxzxzxzzxzzzzzzzxzxzzzzzxxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
