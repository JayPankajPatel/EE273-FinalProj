class c_1043_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1043_6;
    c_1043_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01z00010xzzzxz000x0z0zzxzz1x0z10zxzxzxzxzxzzzzzxxzzxxxzxzxxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
