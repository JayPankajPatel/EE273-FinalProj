class c_1037_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1037_6;
    c_1037_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0zxx1zzx00zxz00z01x00xx0z1x011xxzxxzxxxzzzzxzxxxzzxxzzzzzxxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
