class c_1627_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1627_6;
    c_1627_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z00zzxzx1x11zxzxzz010zxz101xz1x0xxxzxxxxzzxzzxxxzxzzzzzxxxzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
