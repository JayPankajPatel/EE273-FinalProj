class c_1241_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1241_6;
    c_1241_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00z10x1xxxz100x1xxz0101z0x0xxzx0zxxzzxzxxxzxzxzxxxxxxxzxzzzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
