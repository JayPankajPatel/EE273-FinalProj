class c_1657_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1657_6;
    c_1657_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxx11z0x0xzxz01x000x1z1xz11zz01xzzzzzzzxxxxxzxzxzzxxxxxxxxzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
