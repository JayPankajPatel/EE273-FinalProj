class c_1571_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1571_6;
    c_1571_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0z1zzx0zzzz1x1zzz0xx100xzz0zzzzxzzxzzxxzxxzzxzzxzxxxzzzxzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
