class c_126_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_126_6;
    c_126_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zxzzx1100xxzzxxz00zxzzz0x1z0xx0xxxxxxxzzxzzzzxzxxzzxxzzzzzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
