class c_1862_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1862_6;
    c_1862_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzz0011xzz01xzx0x001x101zx1xz11zzxxxzxzzzzxxxzxzzxzzxxxxzxxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
