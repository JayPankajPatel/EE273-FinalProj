class c_40_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_40_6;
    c_40_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxxxx1x0xz001xxz0010zx1xx1zz11xzzzzxxxzxxxxzxzxzzzxxzxxxzzxxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
