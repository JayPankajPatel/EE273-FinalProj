class c_462_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_462_6;
    c_462_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x0000001z00xx0zz1z0z01xz01zxz0xxxzzxxzxzxxxxxxzxxxxxzxxxxxzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
