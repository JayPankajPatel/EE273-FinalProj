class c_1822_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1822_6;
    c_1822_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx010z1xxx11zz01xx0zz00x00100zzxzxxzzxxxzxxzxxzxxzxxxzzzxzzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
