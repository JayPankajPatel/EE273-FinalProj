class c_1747_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1747_6;
    c_1747_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11x10z11z11z10xzx0z1xxxx0x0z0x11zxxzxxzzzxzxzxxxxzzxzzxxzxzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
