class c_521_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_521_6;
    c_521_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1xxxx001x0zxx11100xxz00xxxzz0xxxzxxxzzzxxxxzxxzxzxzzzzzxzxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
