class c_879_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_879_6;
    c_879_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xxz0x10zzx0x1zz1xzzz0zz1zxx0zz0zxzxxzxzxzxzzzxzxxxzzzzzzzzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
