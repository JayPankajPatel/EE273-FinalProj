class c_10_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_10_6;
    c_10_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01xzx11111x10xx01x011zxxx11z1z11zzxxzxzzzxxzxzzzzxzxzxxzzzzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
