class c_1687_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1687_6;
    c_1687_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0100zxxxz100x0z1zx0xxzz1xx1zxzzxzzzxzxzzzzxzzxxxzxzzxxzxzzzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
