class c_1800_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1800_6;
    c_1800_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1xz111z01xz001011x10zz11xz01x11zxxzxxxxxzxxxzzxxxzzzzzxzxzzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
