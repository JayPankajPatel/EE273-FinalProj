class c_790_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_790_6;
    c_790_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x11z0zz10110xz1x00000xz00z101z1xzzzxzzzzxxxxxxxxxxxzzxzzxzxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
