class c_1673_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1673_6;
    c_1673_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z0011z11100zzz100z01x1z00xzzx0zzzzzxzxxzxxzzzzzzxxzxzxzzzzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
