class c_876_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_876_6;
    c_876_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00x0zz0xz011zx0z01xzxzz1z10z1z11zzzxxxzzzzzzxzxxzzxxxzxzxzxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
