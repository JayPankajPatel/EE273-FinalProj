class c_1707_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1707_6;
    c_1707_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01z1z10x101011z0zzzz01zzz0xzzzz1xzzxzzzxzxxxzxzxxzzzzxzzxzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
