class c_1209_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1209_6;
    c_1209_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00z10z1x0zx10zx0zzx1z0z0000xzzx1zzzzxzzxzzzzzzxxxxzzzxzzzxxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
