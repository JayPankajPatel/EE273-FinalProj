class c_809_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_809_6;
    c_809_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x010zzzz001zxzxxx01xxz01xz1z111xxzzxzxxxzzzxxxxzzxxxxzxzxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
