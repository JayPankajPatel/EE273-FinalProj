class c_1777_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1777_6;
    c_1777_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz1zzx1z0z1zzz010zz110x1x0xxx101xxzzxzzzxzxzzxzxxzxxxzzzzzzxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
