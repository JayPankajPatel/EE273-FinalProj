class c_905_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_905_6;
    c_905_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx0000z1x0z0z00z0zzx00x01xz0zx0zxzxzxxxzzzzxxxzzzzxxxzxzxzxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
