class c_1270_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1270_6;
    c_1270_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xx10zz11z0xz01z0zx11zxzzzzx0xz1xzzzzxzxzzzzzxzxxxxxxxzzzxzxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
