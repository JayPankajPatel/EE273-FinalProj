class c_1592_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1592_6;
    c_1592_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z00z1xzx1xx000100x11x1zz00z00z0zzxzzzxzxzxxxxxxzzzzzxxzzzxxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
