class c_72_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_72_6;
    c_72_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01z0110z11z000zz001zx0011xz1x1xxzzxzxxxzzxxzzzzxxxzxxxxxzxzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
