class c_471_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_471_6;
    c_471_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01z1z010x0zx11x0000000z110zz0x01xzzxxxxzxzxxxzxxxzxzxxzxzzzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
