class c_489_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_489_6;
    c_489_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0zxzx1001001z0xzxz1x10x1x1z110zxzzzzxxxzxxxzzzxzzxzzxxxxxxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
