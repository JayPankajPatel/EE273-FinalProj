class c_22_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_22_6;
    c_22_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1xxxx000x1111zzzxxxxx0x0z110z01zzzzzzxxzzxzxzzxxxxzxzxzzzxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
