class c_1723_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1723_6;
    c_1723_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xxz00x0xz0xz1z0xz0z0x0zx0z0z11zxzzzxzzxxzxxzxxxxxzxzxxzzxzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
