class c_1672_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1672_6;
    c_1672_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0x01xxxzxz1xzxz1zz00xxx0100zzx0xxxxzzxxzzzxzzxzzxxxzzzxxxxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
