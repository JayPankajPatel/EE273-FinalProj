class c_1420_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1420_6;
    c_1420_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z01xx0xz1z11zz111z0x1z0zzz000z1xzzzzzxxxzxxxzxxxxzzxzxzxxxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
