class c_1539_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1539_6;
    c_1539_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10000x000001x00010xxz1xzzxz1z0x0zxxzxzxzzxzzzzzxzxxzxxxzzzxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
