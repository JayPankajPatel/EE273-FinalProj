class c_1779_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1779_6;
    c_1779_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0xz0x0zx1zx1z1z0z1zxx000xx10x00zxxxzxxzxxzzzzxxxxzzzzzxxzzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
