class c_1590_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1590_6;
    c_1590_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz0110xzzxx0zz1zz10xxx10zxx1xx1zzzzxzzzxzzzxxzzzzzzzzzxxzxzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
