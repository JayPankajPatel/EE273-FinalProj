class c_1610_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1610_6;
    c_1610_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xx0z1x0x1zz1x1x00zzx110zzzz1xx1zxzzxzxzxzxxzzzzxxzxxzxxzxzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
