class c_1331_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1331_6;
    c_1331_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z10zx0zzx1z1z0010x0xzz00zz11zzxzzxxxzxxzzzzxxzxzzzzzxzzxxzzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
