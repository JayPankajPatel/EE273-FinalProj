class c_253_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_253_6;
    c_253_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10z11zzx1x1xzxzz0zzz1x0xx010x1zxzzzxxxxzxxzzxxxxxzzxzxxzzxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
