class c_1752_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1752_6;
    c_1752_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx1z11zxzx1z10111x1xx0zzxx011xzxxxzzxzzxxzzzzxxxzxzxxzzzxzzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
