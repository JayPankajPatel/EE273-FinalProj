class c_1836_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1836_6;
    c_1836_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zxz0zzz1xx0x000xzzzxx1xxxzx1zz1zzxxzxzzzzzzxzzzzxxzzxzzzxxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
