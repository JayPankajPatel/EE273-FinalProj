class c_1608_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1608_6;
    c_1608_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1000zx0110xxx1011zzx111zxz1z1x0xxzxzzzzzxxxzxzxxxzxxzxxzzxzzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
