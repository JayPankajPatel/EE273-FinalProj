class c_962_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_962_6;
    c_962_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zzxzxx11101x1x11x01011100xx0xx1xxxxzzxxzxxzzxxxxxzzxzxzzxxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
