class c_1712_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1712_6;
    c_1712_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0101010x1010z101zx1xzxzx0z1xzzxzxxzxzzzxxxzzxxxzzxxxzxxzzzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
