class c_275_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_275_6;
    c_275_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00zx1100xz0x0x1x1z11110xxz10010xzxzzzxxzzxzzzzxxzxzxxzzxxzzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
