class c_1427_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1427_6;
    c_1427_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx0x100xz00xxxzx100zxxxxxz0x01x1zxzzxxxzzzzzzxxxxzzzxxxxzxxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
