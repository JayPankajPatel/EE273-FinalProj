class c_371_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_371_6;
    c_371_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz10010zxx1z0x0xxxz10x01xz0z10x1xxxxxzxxzzxzxzxxzxxzxxzzzzzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
