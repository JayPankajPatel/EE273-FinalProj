class c_1833_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1833_6;
    c_1833_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1110zx0x0x10x1xx1x00xz1000zz1x1zzxzzzxzxxzzzzxxxxzzxzzzzzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
