class c_477_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_477_6;
    c_477_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xxz0z111000001x1x00xzxxx1zzzx10zzzzzzzxzzxxzzzzzxxzxzxzxxzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
