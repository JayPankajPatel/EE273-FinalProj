class c_1493_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1493_6;
    c_1493_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0111111x0x0zzzzzz00z0x1x01zxxxzzzxxxxxzzzzxxzxzxxzxxxxzzxxxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
