class c_570_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_570_6;
    c_570_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzzxxzzz011x101x10xz110z0zxxx11zxxzxxxzzxzxxzxzxxxxzzxzxxxxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
