class c_252_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_252_6;
    c_252_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1010zz1z0zxx10zzz000100110xzxxxxxxxxxxzxxxzzzzxxxzxzzxzzzxzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
