class c_1176_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1176_6;
    c_1176_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x100x10zzx0zzzzz11x01zx0x1x10z1zzxzzzzxxxzzzzzxxzxxzxzxxzzxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
