class c_91_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_91_6;
    c_91_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxz110zz0z0x0zz0zz110zx100zz01zxzzzzxzzxxzxxzzzxxzzzzzxxzxxzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
