class c_1289_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1289_6;
    c_1289_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01x0x1xxxx0z0zx00zxxzxz0z010001zxxzxxzzzzxxxzxzxxzzzxxxxzzzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
