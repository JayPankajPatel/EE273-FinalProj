class c_356_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_356_6;
    c_356_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00xz1zx1z1000x00zzx01z0x0x01x0zxxzxxxxzzxzxxzzxxxxzzxxxxzzxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
