class c_1030_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1030_6;
    c_1030_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z101zxz110zxz10xxzz11zxz0x111z1xzzxxzzzxzzzzxzxzxzzzzxzzxzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
