class c_833_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_833_6;
    c_833_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0z1zzxzzx11xx10x0x0x0zz0x1z110zxxxxxxzxzxxxzzxxzzxxxzxxzzzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
