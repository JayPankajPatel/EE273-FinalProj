class c_1280_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1280_6;
    c_1280_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xxzzx10x0zx011z1x10x01zx0x0z01zxzzzzxzzxxzxxzzxxzzxzzxxzxxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
