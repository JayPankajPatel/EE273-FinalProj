class c_1549_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1549_6;
    c_1549_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0z1x10zx1xz1zxzz1zxx1xxz001xzx0zxzxzzzzzzzzzxxzxzxzzzzxxzzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
