class c_426_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_426_6;
    c_426_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10xzx000zx0z0000z01x1011zxxxzxz0zxzxzzxxzxxzzxxzzxxzxzxxxxxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
