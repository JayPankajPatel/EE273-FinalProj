class c_1079_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1079_6;
    c_1079_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "001011xzxxz110xx01000z0zzz01z0z0zzzxzxxxxzzxxxxxzzzxzzxzzzxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
