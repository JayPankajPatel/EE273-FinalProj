class c_1765_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1765_6;
    c_1765_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0110z0x0zxz000zzzz0z001x1xx0x0x1zxzzxzxxzzxxzzxzzxxzzxxxxxxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
