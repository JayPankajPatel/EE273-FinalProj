class c_792_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_792_6;
    c_792_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01xzzxzz1zz10xx1zxx1z10x0xzx1x01xxxzxzzxzzzxxzxzxzxzzzzzxxzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
