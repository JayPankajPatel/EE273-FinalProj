class c_992_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_992_6;
    c_992_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00z10z10010xzx0zz1x1000zxx0xxzx0zxxxzxxxxxxzxzxxxxxzxxzxxzzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
