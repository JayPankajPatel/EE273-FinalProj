class c_829_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_829_6;
    c_829_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x0xzxx0xzz0zx1x11x0xx11xx01x110zxzzxxxxxxzxzxzzzzzzxzzxxxzxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
