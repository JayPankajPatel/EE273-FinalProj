class c_583_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_583_6;
    c_583_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1x10zz1001xzx110x010x1zxx1z101zxzzxxxxxzzxzxxxxxxxzzxxxxxzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
