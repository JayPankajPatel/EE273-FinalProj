class c_1061_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1061_6;
    c_1061_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z1xzx01z01xx11xz001z0z0zzz100z1zzxxzxxxzxxxxzzxxxzxzxzxzzxzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
