class c_1243_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1243_6;
    c_1243_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zxzxz11zzxzxxzzz00zxz1xx0x001xzzxzzzxxzzzzxxzzxzxzzxzzxxxxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
