class c_1483_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1483_6;
    c_1483_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11xx0xx11x000zxz10zz1000x1z0z1xxxzzzzxxxzxxzzxzzzzzxzzzzxxzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
