class c_287_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_287_6;
    c_287_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x0zzz0z0z1x10zz1xxxx11x11zzxx0xxzzzxxxxzzxxzxzzzzzxzxxxxxxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
