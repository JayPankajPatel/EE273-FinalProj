class c_1529_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1529_6;
    c_1529_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "010xxxx00xz1x0xzx1zzz11101011110zzzxzxxxzzzzxzzxzzzzxzzzxxzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
