class c_1828_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1828_6;
    c_1828_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1x0z1100zxzz11z1x1000zx00z1xxz1zzzzxxxzzxxxxxxxxzzxzxzzzxxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
