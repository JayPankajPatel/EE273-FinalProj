class c_581_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_581_6;
    c_581_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x11zz1zxxxxz1z100zxxzx10xx11zzzzxxxzzzzzzxzxxxzzzxxzzxzzxxxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
