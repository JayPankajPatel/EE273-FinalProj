class c_1210_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1210_6;
    c_1210_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxxzz0zzx10z1xx110zzx00x0zzx01zzzxzzxxxzzzxzxxzxzzzzzxxzxxxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
