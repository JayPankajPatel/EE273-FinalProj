class c_1659_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1659_6;
    c_1659_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0x01z11zxx1xxzxz1zz0xx1zzx10x0xxzzzxxzxzzzzzzzxxzxxzzxxzxxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
