class c_705_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_705_6;
    c_705_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x1x11z1x001x10011zzz1100x0101z1zzzzxzzxzxxxxxxzxzzxzxzxzzxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
