class c_1172_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1172_6;
    c_1172_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00x0001z00zx1zx1zzzzz1zx001xzxz0xzzxzzzxzzzzxxxzzxxzxxzxzzzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
