class c_701_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_701_6;
    c_701_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx1x11011z10x1z1z1zz0z1xz1x10zzxzzxxxxzzxzxzxxzzzzzxxzzzxxxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
