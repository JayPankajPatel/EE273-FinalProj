class c_672_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_672_6;
    c_672_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x001110xx110x0x11zxz010xzz011z1zxzxxzxzzzzzzxzxxxzxzzxxzxxxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
