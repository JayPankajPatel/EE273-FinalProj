class c_1169_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1169_6;
    c_1169_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01x00001zz11x001xx0zx1zx110z1x11zxzzxzxzxzzzzzzzzzxxzzzzzzzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
