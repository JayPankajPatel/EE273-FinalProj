class c_98_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_98_6;
    c_98_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z101xx0xxz10xxzxz0011zzxz101xxxzzxzxxzzxxzxxxzxxzxzxzxzxzzxzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
