class c_344_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_344_6;
    c_344_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0101xzz0zz00zzzxxzzxz1x00010z0xxzzzxxzzzxxzxzxxxzxzxzxzxxxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
