class c_1880_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1880_6;
    c_1880_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1xzz1zzxzx11z101zx110z10x0zx1xxxzzzxzzzzxxxzxzxxzxxzzxxzzxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
