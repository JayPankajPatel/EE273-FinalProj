class c_1092_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1092_6;
    c_1092_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01x100zz110z101xzx01xxzz1xxz1z10xzzxxzzzxxxzxxzxxzzxzxxxxzzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
