class c_1222_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1222_6;
    c_1222_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0x1111zzxx00111zx0z01x1x01z011zxzzxzzxzxxxzzxxxzxxzxzzxzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
