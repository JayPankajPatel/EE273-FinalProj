class c_1728_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1728_6;
    c_1728_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01zxzxz1x1x1zx100z1x10x01xxxxzx0xxxxzxxxzxxzxzxxzzxzxxxzxzzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
