class c_1499_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1499_6;
    c_1499_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxz0zx0xxx10z0zz110111z001xxx01xxxxxxzzzxzzxxxzzxxzxzzxzzzzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
