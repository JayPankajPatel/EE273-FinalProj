class c_116_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_116_6;
    c_116_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1zxz0x10xzx0z1x0x11x11x0110zzz1zzzxzzzxzxxzzzzzxxxxxzzxxzzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
