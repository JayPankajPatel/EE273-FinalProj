class c_1116_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1116_6;
    c_1116_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00zxx0zzz0xzz0z11x1x110xxz1x0x11xzxxzxxxxxxxxzxxzzxzzzzxxzzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
