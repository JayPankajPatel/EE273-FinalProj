class c_1390_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1390_6;
    c_1390_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "110z01zx1z111x1z1zzxx1xz101x1z1xxzxxxzxxzxxzxxxzxzxzxxzzxzxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
