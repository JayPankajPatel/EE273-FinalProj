class c_626_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_626_6;
    c_626_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z011xx1x00z0xzz0z1z1x1x000xxz1zzxxzzzxzzxxxxxzxxxxxxzzxxzxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
