class c_1738_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1738_6;
    c_1738_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz1z10z0x101x011x01xz0xxx1xzz110zzzzzzxxxxxzxxxzxzxxzxxxzzzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
