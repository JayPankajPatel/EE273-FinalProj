class c_651_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_651_6;
    c_651_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z11x1100x001zxz111xz1z0x1001zxzxxxzxxzzxxxxzzxzxxxxxzxxxxzzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
