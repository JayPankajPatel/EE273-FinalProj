class c_1309_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1309_6;
    c_1309_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxxz1xz1z0zx10110zz10xx0100zx11xxxxzxzzzzzzxzzzzxxzzxxxzxxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
