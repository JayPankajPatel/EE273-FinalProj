class c_1448_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1448_6;
    c_1448_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzzxx1x10x1x1z1xz0x10011zx1z11zzxzxxxxxzxxxzzxxxzxxxxxxzzxxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
