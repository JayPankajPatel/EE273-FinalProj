class c_1757_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1757_6;
    c_1757_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1xzxx0011zz111z0xx01zz0xxzzx1xzxzxzxzxzzzxxxzxzzzzxxxxxzxzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
