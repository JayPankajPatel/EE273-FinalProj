class c_915_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_915_6;
    c_915_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01z1001zz1110x1z111zx100zx01111zzzxzzzzxxzxzxxzxzzzxzzzxzzxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
