class c_1304_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1304_6;
    c_1304_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0zx10x00z11xx1x1x1zxx0xxz0z000zzxzzxxxxzzxzzxxxxxzzxzxzxzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
