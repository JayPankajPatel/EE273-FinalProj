class c_1605_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1605_6;
    c_1605_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x10x001z100110z0x01010011xx1zzxxxzzxzxxzzxxxxzzxzzzzxxxxzzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
