class c_1250_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1250_6;
    c_1250_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxz1z0x0z0x01z0xx01xx0z00x1x10xzzxzxxzxzxzxzxxzzxxxzzxxzzxzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
