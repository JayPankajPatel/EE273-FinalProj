class c_1302_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1302_6;
    c_1302_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx110xxzxx1z1x1zzx110x010x0x11z0xxzxzzzzxxxzxxzzzzzzxxxxzxzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
