class c_108_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_108_6;
    c_108_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx0zxzxzx1x0x0x0zx0000zxz0z1xx1xxzzxxzzzxzzxzxzzxzxxxxzzzzzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
