class c_1557_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1557_6;
    c_1557_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxzzx01z00z11xx1x0x1101010zx01xzxzzzzzzzxzxxxzxzzxxxzxxzxxxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
