class c_545_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_545_6;
    c_545_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01zz0zxz11zx11zz0zxzzx1xxz0x0x10xxxxzzxxxxzxxzzzxzxxxzzxxzxzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
