class c_1032_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1032_6;
    c_1032_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1x0zz0z0zxxx11z1010zx0xzz110z0xzxxxxxxzzzxzxxzxxxzzxxxxxxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
