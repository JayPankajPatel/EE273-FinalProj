class c_1056_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1056_6;
    c_1056_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zx10z11z1100z0xz0x1z0xx010xxz00zxxzxzxxzxzzxzxxxzxzxxzxxzzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
