class c_1200_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1200_6;
    c_1200_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1xxx01z1xzzx11xxxx0z0000zxx000xxxzxzzzxzzxxzxzzzxxxxxxxxzzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
