class c_1709_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1709_6;
    c_1709_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxxxzz10zz0x1z0xzxzxzxzx0110xz10zzzzzxzzzxzxxxxzzxxzzxxxzxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
