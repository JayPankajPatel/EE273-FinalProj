class c_1430_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1430_6;
    c_1430_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1011xx0x11zzx011xzz010z1xxzx0z0xxxzzzzzzzxxzxxzxzzzzzxzzxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
