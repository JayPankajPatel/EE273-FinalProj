class c_1811_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1811_6;
    c_1811_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxx101xzx01z1x11xz1xxzzxzx11xz00zzxxzzzzzzzzxxzzxzzxxzzxzzzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
