class c_218_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_218_6;
    c_218_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0x00101z0zx001z1001zz1100z1zzzzxxxzxzxzzzzxzzzzzxxxzxzzzzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
