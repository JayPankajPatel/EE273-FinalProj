class c_1864_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1864_6;
    c_1864_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0101z000z0x110010xzz0zx110zzzxzxxzzxzxxxxzxzxxxxxxzzxzxxxxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
