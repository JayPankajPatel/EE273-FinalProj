class c_1101_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1101_6;
    c_1101_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0110x1111zz00zzx1zx1xx11xz0x0x0zxxzxzxzxxzzzzxzzxzxxxzxzxzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
