class c_990_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_990_6;
    c_990_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx0000111z0011011zzz0z00z11xz010zzxxxzxxxxzxxxxxxxxzxxzxzxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
