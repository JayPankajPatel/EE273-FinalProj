class c_1231_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1231_6;
    c_1231_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzz01100z1100zx1z1x001zx0xxzz10zzxzxzzxzzzxxzxzzzzzxzxzzxzxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
