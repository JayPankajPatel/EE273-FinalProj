class c_1049_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1049_6;
    c_1049_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx01zxz0xx0zx01z0zz01zxxzx001xzzxxxxzzzxzxzzxzzxxzxzxxzzzzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
