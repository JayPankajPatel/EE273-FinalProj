class c_540_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_540_6;
    c_540_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0xzx001xxxz10z0111z011z0xxxz1zzxzxxzxzxxxxxzzxxxxxxxxzxzxzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
