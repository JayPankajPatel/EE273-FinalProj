class c_1520_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1520_6;
    c_1520_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x11x1xx1xzzz00011z10z0x1x1xx0001xzzzxzzzxzzzxzzzzxxzzxxzzzxzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
