class c_851_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_851_6;
    c_851_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0100z11zx0z0zxzx10zzzzz101zzxxzxxzxxzzxzzxzxzxxzzxzzzzzzxzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
