class c_985_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_985_6;
    c_985_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx11xxz0x000x1x01x1z1010zxx11zzzxzzxxzzxxzxzxzzxzzxxzxzxxxxzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
