class c_973_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_973_6;
    c_973_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z10xx10x11z11xx1000101zxz1101z0zzxxxxzxxzzzzzxzxxzzxxxzxzzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
