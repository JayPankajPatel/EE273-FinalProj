class c_807_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_807_6;
    c_807_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzx0zz11zx00xzzx111z0xzxx01zx11xzzzzxxzzxxzzzzzzzxxxzzzxzxzxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
