class c_1262_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1262_6;
    c_1262_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1001xx1zx1x1zxz00xx10zzzzx00z0zxxxzzzzzzzxzxxxxxzzxzzzzxzxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
