class c_273_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_273_6;
    c_273_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xzz11zz0xz0zx101z00xx10x0x0x00xxxzzzxzxxzxxzzxzzzxxxzzzxxzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
