class c_1342_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1342_6;
    c_1342_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z11zz01zzxxxxx1x1xx00z1z01111z0zzzxxxxxxxzxzxxzxzzxzxzzzxzxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
