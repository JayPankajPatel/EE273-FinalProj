class c_88_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_88_6;
    c_88_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz01zzx1zx1z1zz000x00zz00000xz0zzzzxzzzxzzzzzzzxxxxxzxxzzxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
