class c_1442_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1442_6;
    c_1442_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1011xx1z100000z01xxzzz01z1xz0x1xxxxzzxxxzzxzzxxxzzxzzxzzzxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
