class c_59_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_59_6;
    c_59_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz01zx110xzzxx1000xx1z101xxz11z0xzzzxzxxxzzxzzxzzzxxzzzxxxxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
