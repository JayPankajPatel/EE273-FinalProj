class c_1729_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1729_6;
    c_1729_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z101xxz0111xz0101xxxz1xxx1x11z1zzzzzxzxxzxxzzzzzzxxzxzzxxxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
