class c_226_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_226_6;
    c_226_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x10x0z1zx0x0xzx1x0z011x1xxxxz0xzzxxzzzxzxxzzzxxxzxzzzzzzzxzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
