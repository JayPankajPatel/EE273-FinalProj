class c_1416_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1416_6;
    c_1416_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z010xzxz0x010xzzx010z111zxzzx0x1zxzzzxxxxzxxzzxxxzxxxzzxzzzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
