class c_1572_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1572_6;
    c_1572_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxx01100xz0xz0z01xzx00zx1011zz00xxzxzzxxxxxzxxzxzzxxzxxxzzzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
