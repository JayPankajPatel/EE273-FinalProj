class c_690_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_690_6;
    c_690_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z101000xxx101z1z0z11z10z10010x1xzzxxxzzxxzxxzzxxzzxzzxxzxxzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
