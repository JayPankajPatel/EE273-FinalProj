class c_538_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_538_6;
    c_538_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00100xx0z000000011x1zx100011z1zzzxzxxxxxxzxzzxxzxzzzxzxzxzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
