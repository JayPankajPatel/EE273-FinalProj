class c_764_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_764_6;
    c_764_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0z0xzzzzzz0z11x100x1zx1x0z0zzzxxxzxzzzzxxxxzxxzzxzxxxzxzxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
