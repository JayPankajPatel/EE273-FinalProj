class c_268_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_268_6;
    c_268_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0xzx11z0x1xzxxz0xxzxxzx111xz1zzzxzxxxxzzzxzxzzzxxxxzzzxzzzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
