class c_1703_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1703_6;
    c_1703_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00zz0zx10xz00z1x0xx1xz0xz1zx1z11xzxzxxzzxxzzxxxxzxxzzxzxxzxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
