class c_427_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_427_6;
    c_427_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0z10x0zz110xx1x0xx0x11z1xzxz0xxxxzxxxzxxzzxzxxzzxxxzxxxzxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
