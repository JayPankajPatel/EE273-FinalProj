class c_555_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_555_6;
    c_555_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z1xzx00xx1zzz00xz110xzx10z0z01zxxzzzxxzxzxxxzzzzzzzzxzxzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
