class c_465_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_465_6;
    c_465_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11100xzzx1zxxx000xxz0x000xx0z0x0xzxzxzzzxzzxzzzzxzzzxxzxzzxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
