class c_38_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_38_6;
    c_38_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zx101x0z1xx0zxzz0z0xz00x111z10xzzzzzzxzxxzxzzxxzxzzxzzxzxzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
