class c_1502_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1502_6;
    c_1502_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0x0xx0zz0xx11xzzz0xx0z0z1xx110zzxxzzzxxxzzzxzzxxxxzxxzxxxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
