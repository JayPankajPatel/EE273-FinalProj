class c_1582_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1582_6;
    c_1582_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0zxxz10xxzz0z10z0x00zz0z1zx101xzzzxzxzxxxxxzzxxzzxxzzzxzzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
