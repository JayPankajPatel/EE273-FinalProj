class c_1422_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1422_6;
    c_1422_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "100x00z00zzz0z0xxx11x1z00010x1z0zxzxxzzxxxzxxxxzzxxxxxxzxxzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
