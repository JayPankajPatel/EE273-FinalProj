class c_1801_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1801_6;
    c_1801_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zx010x1zxx100x1xx1xxz1xxx1z1xx1xzxxxzxzzzxxxzxzzxxzzxzxxzxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
