class c_1321_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1321_6;
    c_1321_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0101zxxzx0xz01z1001zx1010100x1zzzxzzxxxzxzzxzxxzzzxzzzzxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
