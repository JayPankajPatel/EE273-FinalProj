class c_194_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_194_6;
    c_194_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz00zx0xzx0xzz1z0xzz01z0z1z01zzxzxzxzxxzxxxzzzzzxxxxzxxxzxzxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
