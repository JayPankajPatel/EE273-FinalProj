class c_85_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_85_6;
    c_85_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxz0zzx1zxxx111zz00x1001zzzx11xxzxzxxxzxzzzzzzzxzzxzzxzxxxzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
