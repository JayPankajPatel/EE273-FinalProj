class c_1569_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1569_6;
    c_1569_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "010x1x11011zxxxzxx010xz01z10z0z1xxzzxzzxzzxzzzxxzzzxzxzxxzxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
