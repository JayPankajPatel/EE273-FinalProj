class c_1343_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1343_6;
    c_1343_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z0zzx011z0x0110z1z1z10zzz00z000zzzxxxzxzzzzxzxzzzzxxxxxxzzxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
