class c_1875_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1875_6;
    c_1875_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1xx01x0zzxxz0011101zxzz11zzx1xxxzxzxxzzzzzzxxxzzzzxzzxxxzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
