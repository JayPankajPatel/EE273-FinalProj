class c_706_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_706_6;
    c_706_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx10xx0z1xxzzxz0xzxxzxx1xzx0xz1xzxxzzxxxxxxzzxzzxzxxxzxzxxxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
