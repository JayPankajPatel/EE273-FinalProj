class c_1274_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1274_6;
    c_1274_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxx0x000xxzzz1zxzx1010xzz1001xx1zxzzxzzzzzxxxzxzzxxzxzzzzzxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
