class c_1295_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1295_6;
    c_1295_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1100z0xxxx1x0xz0x11z1z0zxxz00100zzxxxxxzxxxzzzzxzzzzzxxxxxzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
