class c_1802_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1802_6;
    c_1802_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10zxx1z0xx11x01zxz0zzx101x1x0x11zxzxzxxzzxxzzzzxxxxzzzxzxzzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
