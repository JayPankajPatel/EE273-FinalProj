class c_1336_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1336_6;
    c_1336_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz11xxz1010zzzzxxzxx1x0000zx10z0zxxxzzzxzzzzzxxzzzzxxzzxxxxzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
