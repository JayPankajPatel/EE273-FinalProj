class c_909_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_909_6;
    c_909_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00xzx1z1zx0x0z1zzxxxz1zxxz00z0xzxxxxzxzxzzzzzzzxzzzxzzzxzxzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
