class c_720_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_720_6;
    c_720_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz10xzx00zzz11zz0xxzz1xxx1xxx101zzxzxzzxxxzzzxxxxxxzzzzzxzzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
