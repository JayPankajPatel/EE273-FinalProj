class c_1734_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1734_6;
    c_1734_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00z0z00zxzz0x0010zzzx0z11zx1011zxxzxxzzxzzxxxxxzzzxzxzxzxzzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
