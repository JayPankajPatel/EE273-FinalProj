class c_1394_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1394_6;
    c_1394_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zxxzz00010zx0011zz11x1zx0z0x01zzxzzxxxzxzxxzxzzzzzxzxxxzxxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
