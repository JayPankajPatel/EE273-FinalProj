class c_823_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_823_6;
    c_823_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0xz0zzx1xzxz1000xx1010x0z01zzzxzzxxzzxzzxzzzzxzzxxzxxzzxzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
