class c_1838_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1838_6;
    c_1838_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxzz0000zxx00011zzxz0xz001x0xz01zxzxxxxxxzxzzzxzzxxzxxxzzzzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
