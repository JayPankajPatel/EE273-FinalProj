class c_1256_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1256_6;
    c_1256_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11z11z0x000000x1101z10zx101x1z10zzzxzzxzzzzxzxxxxxxzzzzzzzzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
