class c_1135_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1135_6;
    c_1135_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx0x00zz0zz1zx00zzxxxx01100x11x0zzzxzzzxzzzzzxxxxzzzzzxzxxzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
