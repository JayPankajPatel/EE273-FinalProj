class c_1369_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1369_6;
    c_1369_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11z1x1zz00z1zz101z0z0z0x0zzxxxx0xxxxzxxzzzxzxxxzzxzzzzzzzxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
