class c_1227_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1227_6;
    c_1227_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzzx000x11zzxzx11x1z000011xxx11zzzxxxzxxxzzxzzxzzxzxzzzzzxxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
