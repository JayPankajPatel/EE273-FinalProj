class c_1795_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1795_6;
    c_1795_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1001zz110z1zzxx1x0xxxxz0x1z0000xxzzxzzxxzxzzxzxzxxzxxxzzxxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
