class c_281_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_281_6;
    c_281_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xx01z1zx001xzxx1x11101z010011xxxzzxzxzxzxxzzxzxzxzzxzxzzzxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
