class c_1360_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1360_6;
    c_1360_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zx10001z1xxx1zz0x0xxzxxz1x011xzxzxxxxxxxzzzzzzzzxzzxzzxxxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
