class c_1553_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1553_6;
    c_1553_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzxxzx11z01x0zx0z011xzzzz010xx10xzzxzxxzxzxzxxxxzxxxzxxxzzxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
