class c_244_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_244_6;
    c_244_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzx0111x0zx000z0z101xx0xz1xzx11xzzxzxxzxxxzzzzzxzxxxxzzxzzzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
