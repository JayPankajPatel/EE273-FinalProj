class c_65_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_65_6;
    c_65_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z0zzz010xx00z00xxzzz0zzzz00z000xzxxzzxxxxxzzxzxxzzxzzxxxzxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
