class c_1715_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1715_6;
    c_1715_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11x0xzz0zzz1101xxx0xzz01110x0x00xzzxxxxxxxxzzzzzzxxzzzzxxzzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
