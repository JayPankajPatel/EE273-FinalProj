class c_1585_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1585_6;
    c_1585_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11x00zzz1xxxz11x0x1xz001x0zxxxz1zzxxzzzzxzxxzxzzxxzxxxzzxzzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
