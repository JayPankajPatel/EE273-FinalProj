class c_818_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_818_6;
    c_818_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z1101xzx0x101zx010z0x1z1z1001xzxxzzzxxzxzxxzzxxzzxzzzzzzxzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
