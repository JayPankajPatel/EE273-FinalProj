class c_1085_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1085_6;
    c_1085_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x01000010x1z0x111111zzzx0x00zzxzzzzzzxxzxzxzxzzxxxzzzxxxxxzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
