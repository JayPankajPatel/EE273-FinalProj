class c_1229_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1229_6;
    c_1229_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx1zz0xx0110001xx0001xz0z01x00z0zzxzxzxzxxzxzxxzxzxxxxxxxxxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
