class c_1181_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1181_6;
    c_1181_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x00zzz11zz11zx10z1x0x10100111x1xxxzzzxzxxxxzzzxzzzzzxxzzxxzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
