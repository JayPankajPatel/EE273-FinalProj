class c_1399_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1399_6;
    c_1399_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0z1000zz110zx00010100x011z01z0zxzzzzxzxxxxxzzxxzxzxzzzxxxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
