class c_1829_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1829_6;
    c_1829_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01zz11101zz00zzx00z100zzz1x0100xxxxxzxxxxzzxzxxzxzzzzzxxzxzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
