class c_9_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_9_6;
    c_9_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xz011z1x10x01zz1z01z1zxx00101xzxxxxzzzxxzzxzxzxzxxzxzzzzxzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
