class c_97_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_97_6;
    c_97_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zxz01zzx01zx1zx11zx010z1x1xzx0xxzxzzzzzzxxxxxzxxxzzxzzzxzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
