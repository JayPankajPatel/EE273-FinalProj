class c_1827_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1827_6;
    c_1827_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z111z0zx100z0z1zzz010xx1zz010x0xxxzzzzzzxxxzxzzxzzzxxzxzzxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
