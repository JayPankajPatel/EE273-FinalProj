class c_1353_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1353_6;
    c_1353_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz10x0x0x0zx1xz1001zzx1z01z1xz0xxzxzzzzzzxxxxxzzzzxxzxxxxzxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
