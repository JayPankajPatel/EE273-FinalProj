class c_1700_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1700_6;
    c_1700_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zz11z01x11x0z01x1110x00x0z110xzzxxxzxzzzxxzxxxxzzxxxzzxxzxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
