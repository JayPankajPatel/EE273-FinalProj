class c_1110_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1110_6;
    c_1110_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z10xx0xxz101xx11x0z1xx0xzzzzz1xzzxzzzzxxzxzzxzxzxzxzzzzzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
