class c_1745_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1745_6;
    c_1745_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz0xxzzz00z1xx1x10100xzzx0zxz011xxzzzzxxxxzzxzzzxxzxxzxzzzzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
