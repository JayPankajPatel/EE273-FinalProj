class c_407_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_407_6;
    c_407_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz10z01zzxx10zz1zx110z00z11x01z0xxzxzzzzzzzxxzzxxxxxzzzxzzzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
