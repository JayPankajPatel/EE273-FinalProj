class c_1746_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1746_6;
    c_1746_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0zxz1x1x0zzxz0zx1zzx0zzz1xxx1xzzxxzxxzxzxxxxzxzxxxxzxzzxxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
