class c_1206_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1206_6;
    c_1206_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00zzzxzzz0xxzzxx1z1x11000xzz1z01xxzxzzzxzzzxzxxzxxxxxxxzzxxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
