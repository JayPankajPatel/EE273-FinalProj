class c_145_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_145_6;
    c_145_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z001zzz00x11z0000x11zzx000z0zzzxxxxzzzzzzxxxzxxzxxzzxxxxzxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
