class c_519_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_519_6;
    c_519_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx01xxz00z1110x10zz0xzxzxxz1zx1xxzzxzxxzxzzzzzxzxxxzzxxxxxzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
