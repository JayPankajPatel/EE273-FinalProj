class c_1775_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1775_6;
    c_1775_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10100xzzz101z1z0x101zxz110xz1x1xzzxxxxxxxxzzxxzxxxzzzzzxxzxzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
