class c_1272_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1272_6;
    c_1272_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xzx01z1x10x0xxx010zz0x1xz0111xzxzxxxzxzzxzxxzzxxzzzxxxzzzxxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
