class c_1472_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1472_6;
    c_1472_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxxx0zz0xxzz0x1x01zz11x1zz1xx00zzzzxxxzxzzxzxxzxxzxzzxxxzzzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
