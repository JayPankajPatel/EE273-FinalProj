class c_1559_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1559_6;
    c_1559_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1z1001zz0zx100xx101xz0z11x0xzz0xxzzxzzxxzxzzzzxxzxxxxxzxxzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
