class c_1396_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1396_6;
    c_1396_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx0xx00zx110z01z11zx0zzzxz01zx1xzzxzzxxxxxzxxzzzxzxzxzxxxzzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
