class c_262_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_262_6;
    c_262_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11z00x110x11xx11010xzzxz1zzzxxz1zzzzxzxxxxxzzzxxzxxzzxzxzxxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
