class c_1263_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1263_6;
    c_1263_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzz011zz0z0z1x111zzx01zx1xzz00zzzxxzxzzzzzxzxxxzzzxzxxzzxxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
