class c_1144_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1144_6;
    c_1144_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1010x0zxx1z001zx0x0zzz0zz0zz1z1xzxxzxzxxzzzzzxzzzxzxxzzxzxxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
