class c_969_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_969_6;
    c_969_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0z1000xz011x0zzx111xzx0000xz0xxzzxxzxxzzxzxxxzxxzxzzxzzxxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
