class c_1818_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1818_6;
    c_1818_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1zxz0zxz0110z1zz1x0x1z001z0zxz1zxxxxxzzxxzxxzxxzxxzzxzxzzzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
