class c_848_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_848_6;
    c_848_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x001x11z1010zx1xzx0xzxx0x1010z1zxxzzxxzxzxxzzxxzzzzzxzxzxxzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
