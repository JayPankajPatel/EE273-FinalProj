class c_1517_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1517_6;
    c_1517_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz0x00zz1x1z11zx110z0x0z011zx100zxzxzxzxzzxzxzzzxzzxxxxzzzzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
