class c_1224_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1224_6;
    c_1224_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01zxz011zz01xzx1z100x001100x0x11zzzzxxxxzzxzzzxxzzxxxzxxxxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
