class c_1355_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1355_6;
    c_1355_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx1zxz11011111x11xxzx1x0xz0z11x1xxxzxxxzzxxzxxzzxzzzxzxzzzzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
