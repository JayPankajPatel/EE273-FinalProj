class c_1294_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1294_6;
    c_1294_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1z0zxx10x1zzxzx0z0x1z0xxx000x00xzzxxxzxxzxxxzzxzzzxxxxzxzzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
