class c_827_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_827_6;
    c_827_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxxx1110110xz10xxxx1z001xxxxz00xxzxzxzzzxzzzzzzzzzzxxxzzzxzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
