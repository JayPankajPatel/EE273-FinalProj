class c_1537_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1537_6;
    c_1537_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1010xxx0z1zz1zz1zzxz0zzzzz11x1z1xxzzxzzzxxxzzxxzzxxzzxzzzxzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
