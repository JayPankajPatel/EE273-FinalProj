class c_1090_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1090_6;
    c_1090_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "000xxx110zxxz1zz01z1xzz10x0xxzxzxxzzzxxzzxxxxxzzxzzxxxzzzzxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
