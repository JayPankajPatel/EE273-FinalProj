class c_1246_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1246_6;
    c_1246_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x0x000zxx0x00xzzxz1xxz101x100x1zxzxzxzxzzxxxzxzxzxxzxzzzxxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
