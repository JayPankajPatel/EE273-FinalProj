class c_734_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_734_6;
    c_734_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x1xz011z01z10zzx010zz11100x1xzzxzzzzxzzzzxxxxxzzzxxxxxzzxxzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
