class c_241_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_241_6;
    c_241_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzxzx1zxzzx1x0x11z1zxzxzx11z11xxxxzzxxzxxzzzxxzxxzxzxzzxxzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
