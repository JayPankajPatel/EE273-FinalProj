class c_1683_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1683_6;
    c_1683_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00zxzx00000xxxx10xzz001100x0z1zxzxzxxzxxzxxxxzxzzxzzzxxxxxxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
