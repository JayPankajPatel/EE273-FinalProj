class c_1349_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1349_6;
    c_1349_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz1x0110z0xx11x1z1zzxx1zz0z10zzxzzxzxxzzxxxzxxxzxxzzzxxzxxzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
