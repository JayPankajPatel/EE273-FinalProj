class c_559_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_559_6;
    c_559_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzxx0xzx10z0xz00zx1101zz0xzzz01xxzzzxxzxxzxxzzzzxxzxzzxzzzxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
