class c_1350_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1350_6;
    c_1350_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xx1z00z0x0xz0zz011z0zzzxz01x10zxxxxzxxxzzxxzxxxzxxxxxxxzzzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
