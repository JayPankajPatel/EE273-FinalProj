class c_224_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_224_6;
    c_224_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x1011zz0z10z1x00101z01x1zx100z0xxxzxxxzzzzxzzzzzzxzxxzzzxzzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
