class c_1440_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1440_6;
    c_1440_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "011zx001xz1x1zzz0x1x0x01x10zxxxxzxzzzzzzxxxzzzzzzzxxzzxzxxzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
