class c_867_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_867_6;
    c_867_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11zx11zx11x00z00xzx00xz00xx1001xxzzxzxxxxzxxzxxzzzzzzxxxxxzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
