class c_90_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_90_6;
    c_90_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z01xz10xzx0xxzzxz1xzzxxzxzx1zxzxzzxxxzxzxxzzzzxzzzxxxzzzxxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
