class c_1547_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1547_6;
    c_1547_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1xzx0xx1z0zx10xzxxx1x10zzz0xxx1xzzzxxxxzzzxxzzxxxxzxxxxzzzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
