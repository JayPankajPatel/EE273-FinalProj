class c_1678_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1678_6;
    c_1678_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzzx111x1xxzxzxzx01x1z010z11zx11xxxzzxzxzzzzxxzzxzzxxzxxzxzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
