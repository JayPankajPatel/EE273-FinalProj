class c_1096_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1096_6;
    c_1096_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111z1x10x0xx10zxz0x01zx1x101z1z0zxxxzxxzxxzzxzxzzxxxxzzxzxxxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
