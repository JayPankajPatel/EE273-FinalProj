class c_1187_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1187_6;
    c_1187_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxz01xzz1010x1x0z0xxz0z1xz001xz1zzzxzzzxxzxzzxzzxzxzxzzzzxxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
