class c_1330_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1330_6;
    c_1330_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1x111x1110x0xxx1xx0zx0x00xx100zzxxzxzxxzxxxzxxxxxxzxxzxzxxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
