class c_557_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_557_6;
    c_557_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz1x11zx10xzzz10z01z1x0xzx1xx100zxxzzzxzzxzzxxxzzxxzxzzxxzxzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
