class c_1041_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1041_6;
    c_1041_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x11xx01z0xzxzx0x1x0xxzx111110z0zzzzxzzzzzxxzzxzzxzxzxzzzzzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
