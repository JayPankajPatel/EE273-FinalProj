class c_1654_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1654_6;
    c_1654_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z0z1x11x00z11010010zxz1zz00z000xxzzxzzxxzxzxzzxzxzzzxzxxzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
