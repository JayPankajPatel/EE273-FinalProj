class c_565_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_565_6;
    c_565_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz1x000z1xx01z00xz10zx0zzzx1xx0zzxzzxzxxzxzxxzxxzxzzxzxxxzxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
