class c_1754_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1754_6;
    c_1754_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzz0zzzzz1x01111xxx00x100z1xz11zzzxxxxxxxxzxzxzxzzxxzzxxxzxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
