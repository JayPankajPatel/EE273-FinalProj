class c_1433_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1433_6;
    c_1433_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x1zxzxx0000zz1z0010z0x010xz0zxzxzxxxxzxzxzxzxxxzzxxxxzxxxxzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
