class c_1368_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1368_6;
    c_1368_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz1100zz100z00x0z100zzzxzz0xx000zzxzxzzzzxxzzxxxxxzxzzzzxxxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
