class c_1044_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1044_6;
    c_1044_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxz0011xxzzx01z011xx1zz1zxzx01xzxzxzzxxxxxzzxzzzzxxxzzzxzzzxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
