class c_1402_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1402_6;
    c_1402_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x0x1011z01x0011z10011xx100001z1zxxzxxxzxxxzxzxzxxxxxzzxxxxzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
