class c_210_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_210_6;
    c_210_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x11z0xx000xz00x101100x11xx110z0xxzxzzxxzxxzzzzzzxzzxzxzxxxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
