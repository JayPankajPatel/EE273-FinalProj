class c_114_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_114_6;
    c_114_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zz1zzx100xz011zx1x00x0x1x11x11zzxzzzxxxzzzxzzzxzxzzzxzxxxzzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
