class c_620_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_620_6;
    c_620_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx0z0zz0xzxzz1zzzx01zzz10x0xz110zzxxxxxxxxxxxxzxzxzxxxxzzxzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
