class c_1118_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1118_6;
    c_1118_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzx111zxz1x1zzx1110z1010x0x11xz0zzzzzzxzzxxxzxzxxzxxzxxxzzxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
