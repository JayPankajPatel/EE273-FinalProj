class c_1560_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1560_6;
    c_1560_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0zxx01x10x011z0zx1z1zx00xzxx0xzxxzzxzxzzzzxxzxxxxxxxxzxzzxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
