class c_1785_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1785_6;
    c_1785_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z11xz001zx10zx01z01zxxz1zxz0xxxxxxzzzxxzxxzxxzzzzzxxzxxzxzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
