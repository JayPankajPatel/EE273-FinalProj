class c_1286_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1286_6;
    c_1286_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzx10xx1xzz111010x1xz1z1101zz11xzzzxzxxxzxzxxxxxxzzzxzzzxxxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
