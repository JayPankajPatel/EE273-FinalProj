class c_951_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_951_6;
    c_951_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01x011xx11x0xxzx100101z00z1zzzx0zzxzzzxzzxxxzxzzxxzzxzxxzzzxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
