class c_1855_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1855_6;
    c_1855_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz010x001x0x0zzxxz0zx0zx11xz11z0xxzxxzxzzxzxzxzzzxxzxxxzzzzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
