class c_1776_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1776_6;
    c_1776_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx0x1zx0zx00x0010100x1zzxxxzx000zxxxxzzxxxxxxzzxzzxzzzxzzzxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
