class c_1587_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1587_6;
    c_1587_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10z000zzx1x0011z10xx0001z001x0xzxxxzzzzxzzzxxxxzzxzzxxzxzzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
