class c_71_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_71_6;
    c_71_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00z00z0z01zx10zxz010zxxxzxx0110xzxzxxxzzxxxxzxzxzzxxxzxzzzxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
