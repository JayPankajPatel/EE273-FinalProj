class c_135_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_135_6;
    c_135_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zzx10x00z1z1xxx00x10z0z1x01z01xxzxzzxzxxzzxxxzxzzxxzzzzxxzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
