class c_79_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_79_6;
    c_79_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1000zz10xx101x01xx1xx0xxz01zxxzxzzzzxzzxxxzxxzzzxxzzxxzzxxzxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
