class c_1358_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1358_6;
    c_1358_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1111xx10x0000zx11xzz1011xxzz0x1xxxzzzzxzxxxxxzxzzzxxzxzzxzxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
