class c_1690_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1690_6;
    c_1690_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1011z1101z0011x0x001xz1100zz1z1xzzzxxzxzxzxzzzxxzzxxxxzzxxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
