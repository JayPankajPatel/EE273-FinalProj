class c_1105_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1105_6;
    c_1105_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x1100zx1zxzx1z1x11z1111x0z111z0xxxzzxzxzzzxzzzzxzzzzzxxxxzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
