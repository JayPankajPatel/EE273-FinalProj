class c_457_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_457_6;
    c_457_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00x0xxz001zxxz110z1zz110010z1z11zzzzxxzzzzzzzzxxxzzzzxzzzxxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
