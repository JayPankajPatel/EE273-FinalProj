class c_1597_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1597_6;
    c_1597_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "101z1001z1z0zzxxx1zzz01x0x000010xxzzzxxzxzxzzzzxxxzzzxxzzxxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
