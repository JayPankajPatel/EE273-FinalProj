class c_107_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_107_6;
    c_107_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "110zzzzx0101z10xz0zx0xz0100z1x0xxzxzxxzxzxxxxxxxzzzxzxxxzzzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
