class c_526_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_526_6;
    c_526_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x101x01zxzxzx011zxz010xz0z10xzzzzzzxxzxxxzxxxxzzxxzxxxxzzzzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
