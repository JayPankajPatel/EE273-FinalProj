class c_136_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_136_6;
    c_136_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zxxz11x0xz010110110000x0001z00xxxzxzxxzzzxxxxzzzxxzxzxxzxxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
