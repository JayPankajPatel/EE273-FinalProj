class c_1327_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1327_6;
    c_1327_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zxz0xz0z0000x00x1xz010zzz0x0zz0xxzxzxzzxxzxzxzzxxxxzxzzxzxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
