class c_1264_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1264_6;
    c_1264_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11z100111zxzx01zzzz1z10101zx0x11zzzxzxxxxxzzxxxzxzzxzxzzxzzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
