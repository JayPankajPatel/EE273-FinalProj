class c_1637_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1637_6;
    c_1637_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0xzxx010x00x0z01xx10xx0zxz0zzx0zzxzxxxxzzxzxzxxzzzzxxzzxzxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
