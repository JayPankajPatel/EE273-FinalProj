class c_81_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_81_6;
    c_81_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x10111z0x01z0xxxzzx1zz101xx1zzxzxzzxzxzzxzxxzxzxxzxxzzxxxxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
