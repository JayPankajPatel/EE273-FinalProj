class c_1237_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1237_6;
    c_1237_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxx111x1x001x011z01z110x000z11xzzzzzxzxzxxxzxzzxxxzzxzxxxzzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
