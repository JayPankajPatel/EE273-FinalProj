class c_820_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_820_6;
    c_820_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z101xx0001x10zz0xz1xx001zxzzx1zzzzzxxzxzxxzxxzzzzxzxxzxzxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
