class c_774_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_774_6;
    c_774_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0101100zxzxz10zxzxxxzx1zz11xxzxzxzxxzxzzzxxzzxxzzxzxzxxzxxzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
