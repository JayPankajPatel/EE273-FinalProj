class c_11_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_11_6;
    c_11_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10xzxz10x001xz0x001100z10x01z0zxxxzzzzxxzzxxxzxzzzzxzxzzzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
