class c_884_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_884_6;
    c_884_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xxz011xzx11xx0zz11zzzz0z1xx0zz0xzzxzzzxzxzzxxxzxzzxxxxzzxzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
