class c_1486_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1486_6;
    c_1486_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0z0000zzz0xxxz0z0z1xx0xxzzz000zxxxzzzxxxxxxxxxxxzxxzzzxzxzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
