class c_604_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_604_6;
    c_604_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xzxz10zzx0zxzxx0x1xxx1xx10x0xx1zzzxzzzxzxxxzxxxxzxxzxxxxzzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
