class c_389_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_389_6;
    c_389_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z01zxzzzzz110zx0z000z001x110xxxxxxxzxxxxzzxxxxzzzzxxxzzzxxzxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
