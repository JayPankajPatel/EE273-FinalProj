class c_1051_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1051_6;
    c_1051_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zz0zzxx00z1xx0z1z01x0xxz10zzz0xzxxzzzxzzxzzzxxxxxxzxxzxxzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
