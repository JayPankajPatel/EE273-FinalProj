class c_717_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_717_6;
    c_717_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00001zzx00xx11z0xzzz1zz0z0z1001zxzxxzzzzxxxzxzxxzxzxxzxxxzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
