class c_1858_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1858_6;
    c_1858_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x00xx0z10zz0zx1001z111110x0x001zxxxxxxzzzzxzzxzxxzxzzzzzzzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
