class c_1600_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1600_6;
    c_1600_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1000xxz0x101x000100z0z01xx10z1zxzxzzxxxxxxzzxzxzzxxxzzxzzxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
