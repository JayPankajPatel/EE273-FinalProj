class c_1400_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1400_6;
    c_1400_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xz100110zx00z000010xzxx0x10z00xxzxxxzzxxzzxzxzxzxzxzxzzzzxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
