class c_1357_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1357_6;
    c_1357_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x0zxxxzxxx1z0z111x000zx01x100x0zzzzzxzxzzxzxzxzxzxxxzxxzzzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
