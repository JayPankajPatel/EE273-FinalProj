class c_113_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_113_6;
    c_113_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1xz1zx00110x11xxx0xxxx0xz0x010zzxzzxxzzxxzxzzxzzxzzxzxxzzxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
