class c_1292_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1292_6;
    c_1292_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0z0z11x0xxxzz0xxx011101zxx0xxz1zzxzxxxxzzzzxxzzzxxxzxxxxxzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
