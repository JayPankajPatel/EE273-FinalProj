class c_1848_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1848_6;
    c_1848_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x0xzzzx00zxzzz1011xxz11xxz001z1zxzzxxzxxzxzxzzxzzzxzzxxxzzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
