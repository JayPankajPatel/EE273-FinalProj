class c_702_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_702_6;
    c_702_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111xz111zxx1zz010x0011x000xz1z1zxzxzxzzxzzzxxxzzzzzxzzxxzxxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
