class c_1684_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1684_6;
    c_1684_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11xz0z1x0x1xxx0101xxzz0z101zxzx1zzzzzzzxxxxxxxxxzxzxzzxxxxzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
