class c_1469_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1469_6;
    c_1469_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxz011x1101zz01011x1z1xxx1xx10xxzxzzxzxxxxzzxzxzxxzxxxxxxxzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
