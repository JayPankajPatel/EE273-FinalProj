class c_1562_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1562_6;
    c_1562_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxx1x0x0x0z001z1zz00x1zx010z11xzxxxzzzzzzzxzxzxxzzxzzxxxzzzzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
