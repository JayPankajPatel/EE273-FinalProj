class c_12_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_12_6;
    c_12_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01x1x0xzzzx11z1z1xxx10x1x1x0101zzxxxzxzxzxzzxzzzxxzzxxzzzzzxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
