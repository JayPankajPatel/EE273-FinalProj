class c_712_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_712_6;
    c_712_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10000z000zz0zzz1xz0z1z01x1x0010zzxxxzxxxzxxxxzxxxzzxxzzzzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
