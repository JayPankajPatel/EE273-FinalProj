class c_573_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_573_6;
    c_573_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x1z0x0xxx1x0x010011xxzx01z0x111xzxzxzxxzzxzzxxzzxzxzxxzzxzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
