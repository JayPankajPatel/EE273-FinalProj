class c_1883_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1883_6;
    c_1883_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0zxzz0x0zzz0111xx1z0111x1z0xzzxxzxzzzzxxzzzzxxzzzxzzzzxxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
