class c_70_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_70_6;
    c_70_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0zz0zz1110zz010011zzz1001z11z1zzzxxxzxzxzzxxzxxxxxxzxzxzzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
