class c_58_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_58_6;
    c_58_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z111z01zxz110x111x1zz1zx10x0zzxxxxzxzxzzzzzzxxzxxzzxxxzxxzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
