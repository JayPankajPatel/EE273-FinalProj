class c_830_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_830_6;
    c_830_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzx0x11xz00100x0zx1z00xz01xx11zxxxzxzzzxxxzzxzxzzxxzzxzzxzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
