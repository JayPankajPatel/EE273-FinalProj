class c_1589_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1589_6;
    c_1589_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1xx11zxzxzz1z1zz0z0x00zx11z101xzxxxzxzxzxxzxzxzzzxzzzxzzzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
