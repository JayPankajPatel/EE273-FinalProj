class c_251_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_251_6;
    c_251_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz0zzzxzxz0010x0x0x100z1x0100xzzxzxxzzxxxzzzxzzzxzzzxzxxzxxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
