class c_1162_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1162_6;
    c_1162_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zx000xxxxx0011xxz0z010x1xx0x11xxzxzxzxxxzzzxzxxxxxzxzxxxzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
