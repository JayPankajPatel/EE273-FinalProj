class c_27_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_27_6;
    c_27_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z00x1xz00x0z10xxz1zzz011z10zx0z0zxxxxzzxxzxzxzzzxzzxzzzzzxxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
