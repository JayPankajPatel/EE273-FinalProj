class c_901_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_901_6;
    c_901_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zx11zz1zz0x10zx111z110z00z0x01zzxzzxzzxxzxzxzxxzxzzxzxxxzzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
