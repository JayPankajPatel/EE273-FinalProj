class c_1120_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1120_6;
    c_1120_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "110zzzz1z0xx0zxzz1z1zzx1xzzzxxzxxxxxxzxxxxxxzzxxzxxxxxzxxzxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
