class c_822_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_822_6;
    c_822_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x1x011xx00x1xxz10z1xx00x10111z0xxxxzzxxxzxzzzzzzxzxxzzxxzzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
