class c_546_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_546_6;
    c_546_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zxz1xz0zxx001110zzxxzx11z0xxz01xxzxzzzxzzzxxzzzzxxxxzxzxxzzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
