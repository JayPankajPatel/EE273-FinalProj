class c_1257_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1257_6;
    c_1257_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xxz1zz0z00z0x1zzz1xz00zz000x11xxxxzzxzzxzxzxxxxzzxxzzzxxxzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
