class c_358_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_358_6;
    c_358_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z00xx11zz0xz11zxxz10x00zzxx11x1zzzzxzxxxxzxxxzzzzxzzzzxxzzxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
