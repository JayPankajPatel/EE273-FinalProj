class c_1484_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1484_6;
    c_1484_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz0zzxxz0zx0xz100xxz011xxxzxx011zxxzxxxzxxxxzxzxzzzzzzxzxxxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
