class c_105_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:63)
    {
       (sda_result == 1'h1);
    }
endclass

program p_105_6;
    c_105_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x01zxz0x1xx110000x11zzzz1z01xzzxzxxxzxzzxxxxzzzzzzxzzxzxxxzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
