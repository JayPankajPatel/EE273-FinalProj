class c_1042_6;
    bit[0:0] sda_result = 1'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../seq/tr_paul_sequence.svh:89)
    {
       (sda_result == 1'h1);
    }
endclass

program p_1042_6;
    c_1042_6 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx11x1x0zzxzx1x01z0x0x1zzzz0zx1xzxzxzxzxxxzxxxxxxxzzzxzxxzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
